`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Lena Voytek
// 
// Create Date: 11/22/2018 03:32:35 PM
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top(Clk, MemAddress, WindowAddress, MemWrite, MemRead, WriteData, SAD_out );

    input Clk, MemWrite, MemRead;
    input [31:0] MemAddress, WindowAddress, WriteData;
    
    output wire [31:0] SAD_out;
    
    wire [31:0] AD0_in_A,
                AD0_in_B,
                AD1_in_A,
                AD1_in_B,
                AD2_in_A,
                AD2_in_B,
                AD3_in_A,
                AD3_in_B,
                AD4_in_A,
                AD4_in_B,
                AD5_in_A,
                AD5_in_B,
                AD6_in_A,
                AD6_in_B,
                AD7_in_A,
                AD7_in_B,
                AD8_in_A,
                AD8_in_B,
                AD9_in_A,
                AD9_in_B,
                AD10_in_A,
                AD10_in_B,
                AD11_in_A,
                AD11_in_B,
                AD12_in_A,
                AD12_in_B,
                AD13_in_A,
                AD13_in_B,
                AD14_in_A,
                AD14_in_B,
                AD15_in_A,
                AD15_in_B,
                AD16_in_A,
                AD16_in_B,
                AD17_in_A,
                AD17_in_B,
                AD18_in_A,
                AD18_in_B,
                AD19_in_A,
                AD19_in_B,
                AD20_in_A,
                AD20_in_B,
                AD21_in_A,
                AD21_in_B,
                AD22_in_A,
                AD22_in_B,
                AD23_in_A,
                AD23_in_B,
                AD24_in_A,
                AD24_in_B,
                AD25_in_A,
                AD25_in_B,
                AD26_in_A,
                AD26_in_B,
                AD27_in_A,
                AD27_in_B,
                AD28_in_A,
                AD28_in_B,
                AD29_in_A,
                AD29_in_B,
                AD30_in_A,
                AD30_in_B,
                AD31_in_A,
                AD31_in_B,
                AD32_in_A,
                AD32_in_B,
                AD33_in_A,
                AD33_in_B,
                AD34_in_A,
                AD34_in_B,
                AD35_in_A,
                AD35_in_B,
                AD36_in_A,
                AD36_in_B,
                AD37_in_A,
                AD37_in_B,
                AD38_in_A,
                AD38_in_B,
                AD39_in_A,
                AD39_in_B,
                AD40_in_A,
                AD40_in_B,
                AD41_in_A,
                AD41_in_B,
                AD42_in_A,
                AD42_in_B,
                AD43_in_A,
                AD43_in_B,
                AD44_in_A,
                AD44_in_B,
                AD45_in_A,
                AD45_in_B,
                AD46_in_A,
                AD46_in_B,
                AD47_in_A,
                AD47_in_B,
                AD48_in_A,
                AD48_in_B,
                AD49_in_A,
                AD49_in_B,
                AD50_in_A,
                AD50_in_B,
                AD51_in_A,
                AD51_in_B,
                AD52_in_A,
                AD52_in_B,
                AD53_in_A,
                AD53_in_B,
                AD54_in_A,
                AD54_in_B,
                AD55_in_A,
                AD55_in_B,
                AD56_in_A,
                AD56_in_B,
                AD57_in_A,
                AD57_in_B,
                AD58_in_A,
                AD58_in_B,
                AD59_in_A,
                AD59_in_B,
                AD60_in_A,
                AD60_in_B,
                AD61_in_A,
                AD61_in_B,
                AD62_in_A,
                AD62_in_B,
                AD63_in_A,
                AD63_in_B,
                AD64_in_A,
                AD64_in_B,
                AD65_in_A,
                AD65_in_B,
                AD66_in_A,
                AD66_in_B,
                AD67_in_A,
                AD67_in_B,
                AD68_in_A,
                AD68_in_B,
                AD69_in_A,
                AD69_in_B,
                AD70_in_A,
                AD70_in_B,
                AD71_in_A,
                AD71_in_B,
                AD72_in_A,
                AD72_in_B,
                AD73_in_A,
                AD73_in_B,
                AD74_in_A,
                AD74_in_B,
                AD75_in_A,
                AD75_in_B,
                AD76_in_A,
                AD76_in_B,
                AD77_in_A,
                AD77_in_B,
                AD78_in_A,
                AD78_in_B,
                AD79_in_A,
                AD79_in_B,
                AD80_in_A,
                AD80_in_B,
                AD81_in_A,
                AD81_in_B,
                AD82_in_A,
                AD82_in_B,
                AD83_in_A,
                AD83_in_B,
                AD84_in_A,
                AD84_in_B,
                AD85_in_A,
                AD85_in_B,
                AD86_in_A,
                AD86_in_B,
                AD87_in_A,
                AD87_in_B,
                AD88_in_A,
                AD88_in_B,
                AD89_in_A,
                AD89_in_B,
                AD90_in_A,
                AD90_in_B,
                AD91_in_A,
                AD91_in_B,
                AD92_in_A,
                AD92_in_B,
                AD93_in_A,
                AD93_in_B,
                AD94_in_A,
                AD94_in_B,
                AD95_in_A,
                AD95_in_B,
                AD96_in_A,
                AD96_in_B,
                AD97_in_A,
                AD97_in_B,
                AD98_in_A,
                AD98_in_B,
                AD99_in_A,
                AD99_in_B,
                AD100_in_A,
                AD100_in_B,
                AD101_in_A,
                AD101_in_B,
                AD102_in_A,
                AD102_in_B,
                AD103_in_A,
                AD103_in_B,
                AD104_in_A,
                AD104_in_B,
                AD105_in_A,
                AD105_in_B,
                AD106_in_A,
                AD106_in_B,
                AD107_in_A,
                AD107_in_B,
                AD108_in_A,
                AD108_in_B,
                AD109_in_A,
                AD109_in_B,
                AD110_in_A,
                AD110_in_B,
                AD111_in_A,
                AD111_in_B,
                AD112_in_A,
                AD112_in_B,
                AD113_in_A,
                AD113_in_B,
                AD114_in_A,
                AD114_in_B,
                AD115_in_A,
                AD115_in_B,
                AD116_in_A,
                AD116_in_B,
                AD117_in_A,
                AD117_in_B,
                AD118_in_A,
                AD118_in_B,
                AD119_in_A,
                AD119_in_B,
                AD120_in_A,
                AD120_in_B,
                AD121_in_A,
                AD121_in_B,
                AD122_in_A,
                AD122_in_B,
                AD123_in_A,
                AD123_in_B,
                AD124_in_A,
                AD124_in_B,
                AD125_in_A,
                AD125_in_B,
                AD126_in_A,
                AD126_in_B,
                AD127_in_A,
                AD127_in_B,
                AD128_in_A,
                AD128_in_B,
                AD129_in_A,
                AD129_in_B,
                AD130_in_A,
                AD130_in_B,
                AD131_in_A,
                AD131_in_B,
                AD132_in_A,
                AD132_in_B,
                AD133_in_A,
                AD133_in_B,
                AD134_in_A,
                AD134_in_B,
                AD135_in_A,
                AD135_in_B,
                AD136_in_A,
                AD136_in_B,
                AD137_in_A,
                AD137_in_B,
                AD138_in_A,
                AD138_in_B,
                AD139_in_A,
                AD139_in_B,
                AD140_in_A,
                AD140_in_B,
                AD141_in_A,
                AD141_in_B,
                AD142_in_A,
                AD142_in_B,
                AD143_in_A,
                AD143_in_B,
                AD144_in_A,
                AD144_in_B,
                AD145_in_A,
                AD145_in_B,
                AD146_in_A,
                AD146_in_B,
                AD147_in_A,
                AD147_in_B,
                AD148_in_A,
                AD148_in_B,
                AD149_in_A,
                AD149_in_B,
                AD150_in_A,
                AD150_in_B,
                AD151_in_A,
                AD151_in_B,
                AD152_in_A,
                AD152_in_B,
                AD153_in_A,
                AD153_in_B,
                AD154_in_A,
                AD154_in_B,
                AD155_in_A,
                AD155_in_B,
                AD156_in_A,
                AD156_in_B,
                AD157_in_A,
                AD157_in_B,
                AD158_in_A,
                AD158_in_B,
                AD159_in_A,
                AD159_in_B,
                AD160_in_A,
                AD160_in_B,
                AD161_in_A,
                AD161_in_B,
                AD162_in_A,
                AD162_in_B,
                AD163_in_A,
                AD163_in_B,
                AD164_in_A,
                AD164_in_B,
                AD165_in_A,
                AD165_in_B,
                AD166_in_A,
                AD166_in_B,
                AD167_in_A,
                AD167_in_B,
                AD168_in_A,
                AD168_in_B,
                AD169_in_A,
                AD169_in_B,
                AD170_in_A,
                AD170_in_B,
                AD171_in_A,
                AD171_in_B,
                AD172_in_A,
                AD172_in_B,
                AD173_in_A,
                AD173_in_B,
                AD174_in_A,
                AD174_in_B,
                AD175_in_A,
                AD175_in_B,
                AD176_in_A,
                AD176_in_B,
                AD177_in_A,
                AD177_in_B,
                AD178_in_A,
                AD178_in_B,
                AD179_in_A,
                AD179_in_B,
                AD180_in_A,
                AD180_in_B,
                AD181_in_A,
                AD181_in_B,
                AD182_in_A,
                AD182_in_B,
                AD183_in_A,
                AD183_in_B,
                AD184_in_A,
                AD184_in_B,
                AD185_in_A,
                AD185_in_B,
                AD186_in_A,
                AD186_in_B,
                AD187_in_A,
                AD187_in_B,
                AD188_in_A,
                AD188_in_B,
                AD189_in_A,
                AD189_in_B,
                AD190_in_A,
                AD190_in_B,
                AD191_in_A,
                AD191_in_B,
                AD192_in_A,
                AD192_in_B,
                AD193_in_A,
                AD193_in_B,
                AD194_in_A,
                AD194_in_B,
                AD195_in_A,
                AD195_in_B,
                AD196_in_A,
                AD196_in_B,
                AD197_in_A,
                AD197_in_B,
                AD198_in_A,
                AD198_in_B,
                AD199_in_A,
                AD199_in_B,
                AD200_in_A,
                AD200_in_B,
                AD201_in_A,
                AD201_in_B,
                AD202_in_A,
                AD202_in_B,
                AD203_in_A,
                AD203_in_B,
                AD204_in_A,
                AD204_in_B,
                AD205_in_A,
                AD205_in_B,
                AD206_in_A,
                AD206_in_B,
                AD207_in_A,
                AD207_in_B,
                AD208_in_A,
                AD208_in_B,
                AD209_in_A,
                AD209_in_B,
                AD210_in_A,
                AD210_in_B,
                AD211_in_A,
                AD211_in_B,
                AD212_in_A,
                AD212_in_B,
                AD213_in_A,
                AD213_in_B,
                AD214_in_A,
                AD214_in_B,
                AD215_in_A,
                AD215_in_B,
                AD216_in_A,
                AD216_in_B,
                AD217_in_A,
                AD217_in_B,
                AD218_in_A,
                AD218_in_B,
                AD219_in_A,
                AD219_in_B,
                AD220_in_A,
                AD220_in_B,
                AD221_in_A,
                AD221_in_B,
                AD222_in_A,
                AD222_in_B,
                AD223_in_A,
                AD223_in_B,
                AD224_in_A,
                AD224_in_B,
                AD225_in_A,
                AD225_in_B,
                AD226_in_A,
                AD226_in_B,
                AD227_in_A,
                AD227_in_B,
                AD228_in_A,
                AD228_in_B,
                AD229_in_A,
                AD229_in_B,
                AD230_in_A,
                AD230_in_B,
                AD231_in_A,
                AD231_in_B,
                AD232_in_A,
                AD232_in_B,
                AD233_in_A,
                AD233_in_B,
                AD234_in_A,
                AD234_in_B,
                AD235_in_A,
                AD235_in_B,
                AD236_in_A,
                AD236_in_B,
                AD237_in_A,
                AD237_in_B,
                AD238_in_A,
                AD238_in_B,
                AD239_in_A,
                AD239_in_B,
                AD240_in_A,
                AD240_in_B,
                AD241_in_A,
                AD241_in_B,
                AD242_in_A,
                AD242_in_B,
                AD243_in_A,
                AD243_in_B,
                AD244_in_A,
                AD244_in_B,
                AD245_in_A,
                AD245_in_B,
                AD246_in_A,
                AD246_in_B,
                AD247_in_A,
                AD247_in_B,
                AD248_in_A,
                AD248_in_B,
                AD249_in_A,
                AD249_in_B,
                AD250_in_A,
                AD250_in_B,
                AD251_in_A,
                AD251_in_B,
                AD252_in_A,
                AD252_in_B,
                AD253_in_A,
                AD253_in_B,
                AD254_in_A,
                AD254_in_B,
                AD255_in_A,
                AD255_in_B,
                Adder128_0_in_A,
                Adder128_0_in_B,
                Adder128_1_in_A,
                Adder128_1_in_B,
                Adder128_2_in_A,
                Adder128_2_in_B,
                Adder128_3_in_A,
                Adder128_3_in_B,
                Adder128_4_in_A,
                Adder128_4_in_B,
                Adder128_5_in_A,
                Adder128_5_in_B,
                Adder128_6_in_A,
                Adder128_6_in_B,
                Adder128_7_in_A,
                Adder128_7_in_B,
                Adder128_8_in_A,
                Adder128_8_in_B,
                Adder128_9_in_A,
                Adder128_9_in_B,
                Adder128_10_in_A,
                Adder128_10_in_B,
                Adder128_11_in_A,
                Adder128_11_in_B,
                Adder128_12_in_A,
                Adder128_12_in_B,
                Adder128_13_in_A,
                Adder128_13_in_B,
                Adder128_14_in_A,
                Adder128_14_in_B,
                Adder128_15_in_A,
                Adder128_15_in_B,
                Adder128_16_in_A,
                Adder128_16_in_B,
                Adder128_17_in_A,
                Adder128_17_in_B,
                Adder128_18_in_A,
                Adder128_18_in_B,
                Adder128_19_in_A,
                Adder128_19_in_B,
                Adder128_20_in_A,
                Adder128_20_in_B,
                Adder128_21_in_A,
                Adder128_21_in_B,
                Adder128_22_in_A,
                Adder128_22_in_B,
                Adder128_23_in_A,
                Adder128_23_in_B,
                Adder128_24_in_A,
                Adder128_24_in_B,
                Adder128_25_in_A,
                Adder128_25_in_B,
                Adder128_26_in_A,
                Adder128_26_in_B,
                Adder128_27_in_A,
                Adder128_27_in_B,
                Adder128_28_in_A,
                Adder128_28_in_B,
                Adder128_29_in_A,
                Adder128_29_in_B,
                Adder128_30_in_A,
                Adder128_30_in_B,
                Adder128_31_in_A,
                Adder128_31_in_B,
                Adder128_32_in_A,
                Adder128_32_in_B,
                Adder128_33_in_A,
                Adder128_33_in_B,
                Adder128_34_in_A,
                Adder128_34_in_B,
                Adder128_35_in_A,
                Adder128_35_in_B,
                Adder128_36_in_A,
                Adder128_36_in_B,
                Adder128_37_in_A,
                Adder128_37_in_B,
                Adder128_38_in_A,
                Adder128_38_in_B,
                Adder128_39_in_A,
                Adder128_39_in_B,
                Adder128_40_in_A,
                Adder128_40_in_B,
                Adder128_41_in_A,
                Adder128_41_in_B,
                Adder128_42_in_A,
                Adder128_42_in_B,
                Adder128_43_in_A,
                Adder128_43_in_B,
                Adder128_44_in_A,
                Adder128_44_in_B,
                Adder128_45_in_A,
                Adder128_45_in_B,
                Adder128_46_in_A,
                Adder128_46_in_B,
                Adder128_47_in_A,
                Adder128_47_in_B,
                Adder128_48_in_A,
                Adder128_48_in_B,
                Adder128_49_in_A,
                Adder128_49_in_B,
                Adder128_50_in_A,
                Adder128_50_in_B,
                Adder128_51_in_A,
                Adder128_51_in_B,
                Adder128_52_in_A,
                Adder128_52_in_B,
                Adder128_53_in_A,
                Adder128_53_in_B,
                Adder128_54_in_A,
                Adder128_54_in_B,
                Adder128_55_in_A,
                Adder128_55_in_B,
                Adder128_56_in_A,
                Adder128_56_in_B,
                Adder128_57_in_A,
                Adder128_57_in_B,
                Adder128_58_in_A,
                Adder128_58_in_B,
                Adder128_59_in_A,
                Adder128_59_in_B,
                Adder128_60_in_A,
                Adder128_60_in_B,
                Adder128_61_in_A,
                Adder128_61_in_B,
                Adder128_62_in_A,
                Adder128_62_in_B,
                Adder128_63_in_A,
                Adder128_63_in_B,
                Adder128_64_in_A,
                Adder128_64_in_B,
                Adder128_65_in_A,
                Adder128_65_in_B,
                Adder128_66_in_A,
                Adder128_66_in_B,
                Adder128_67_in_A,
                Adder128_67_in_B,
                Adder128_68_in_A,
                Adder128_68_in_B,
                Adder128_69_in_A,
                Adder128_69_in_B,
                Adder128_70_in_A,
                Adder128_70_in_B,
                Adder128_71_in_A,
                Adder128_71_in_B,
                Adder128_72_in_A,
                Adder128_72_in_B,
                Adder128_73_in_A,
                Adder128_73_in_B,
                Adder128_74_in_A,
                Adder128_74_in_B,
                Adder128_75_in_A,
                Adder128_75_in_B,
                Adder128_76_in_A,
                Adder128_76_in_B,
                Adder128_77_in_A,
                Adder128_77_in_B,
                Adder128_78_in_A,
                Adder128_78_in_B,
                Adder128_79_in_A,
                Adder128_79_in_B,
                Adder128_80_in_A,
                Adder128_80_in_B,
                Adder128_81_in_A,
                Adder128_81_in_B,
                Adder128_82_in_A,
                Adder128_82_in_B,
                Adder128_83_in_A,
                Adder128_83_in_B,
                Adder128_84_in_A,
                Adder128_84_in_B,
                Adder128_85_in_A,
                Adder128_85_in_B,
                Adder128_86_in_A,
                Adder128_86_in_B,
                Adder128_87_in_A,
                Adder128_87_in_B,
                Adder128_88_in_A,
                Adder128_88_in_B,
                Adder128_89_in_A,
                Adder128_89_in_B,
                Adder128_90_in_A,
                Adder128_90_in_B,
                Adder128_91_in_A,
                Adder128_91_in_B,
                Adder128_92_in_A,
                Adder128_92_in_B,
                Adder128_93_in_A,
                Adder128_93_in_B,
                Adder128_94_in_A,
                Adder128_94_in_B,
                Adder128_95_in_A,
                Adder128_95_in_B,
                Adder128_96_in_A,
                Adder128_96_in_B,
                Adder128_97_in_A,
                Adder128_97_in_B,
                Adder128_98_in_A,
                Adder128_98_in_B,
                Adder128_99_in_A,
                Adder128_99_in_B,
                Adder128_100_in_A,
                Adder128_100_in_B,
                Adder128_101_in_A,
                Adder128_101_in_B,
                Adder128_102_in_A,
                Adder128_102_in_B,
                Adder128_103_in_A,
                Adder128_103_in_B,
                Adder128_104_in_A,
                Adder128_104_in_B,
                Adder128_105_in_A,
                Adder128_105_in_B,
                Adder128_106_in_A,
                Adder128_106_in_B,
                Adder128_107_in_A,
                Adder128_107_in_B,
                Adder128_108_in_A,
                Adder128_108_in_B,
                Adder128_109_in_A,
                Adder128_109_in_B,
                Adder128_110_in_A,
                Adder128_110_in_B,
                Adder128_111_in_A,
                Adder128_111_in_B,
                Adder128_112_in_A,
                Adder128_112_in_B,
                Adder128_113_in_A,
                Adder128_113_in_B,
                Adder128_114_in_A,
                Adder128_114_in_B,
                Adder128_115_in_A,
                Adder128_115_in_B,
                Adder128_116_in_A,
                Adder128_116_in_B,
                Adder128_117_in_A,
                Adder128_117_in_B,
                Adder128_118_in_A,
                Adder128_118_in_B,
                Adder128_119_in_A,
                Adder128_119_in_B,
                Adder128_120_in_A,
                Adder128_120_in_B,
                Adder128_121_in_A,
                Adder128_121_in_B,
                Adder128_122_in_A,
                Adder128_122_in_B,
                Adder128_123_in_A,
                Adder128_123_in_B,
                Adder128_124_in_A,
                Adder128_124_in_B,
                Adder128_125_in_A,
                Adder128_125_in_B,
                Adder128_126_in_A,
                Adder128_126_in_B,
                Adder128_127_in_A,
                Adder128_127_in_B,
                Adder64_0_in_A,
                Adder64_0_in_B,
                Adder64_1_in_A,
                Adder64_1_in_B,
                Adder64_2_in_A,
                Adder64_2_in_B,
                Adder64_3_in_A,
                Adder64_3_in_B,
                Adder64_4_in_A,
                Adder64_4_in_B,
                Adder64_5_in_A,
                Adder64_5_in_B,
                Adder64_6_in_A,
                Adder64_6_in_B,
                Adder64_7_in_A,
                Adder64_7_in_B,
                Adder64_8_in_A,
                Adder64_8_in_B,
                Adder64_9_in_A,
                Adder64_9_in_B,
                Adder64_10_in_A,
                Adder64_10_in_B,
                Adder64_11_in_A,
                Adder64_11_in_B,
                Adder64_12_in_A,
                Adder64_12_in_B,
                Adder64_13_in_A,
                Adder64_13_in_B,
                Adder64_14_in_A,
                Adder64_14_in_B,
                Adder64_15_in_A,
                Adder64_15_in_B,
                Adder64_16_in_A,
                Adder64_16_in_B,
                Adder64_17_in_A,
                Adder64_17_in_B,
                Adder64_18_in_A,
                Adder64_18_in_B,
                Adder64_19_in_A,
                Adder64_19_in_B,
                Adder64_20_in_A,
                Adder64_20_in_B,
                Adder64_21_in_A,
                Adder64_21_in_B,
                Adder64_22_in_A,
                Adder64_22_in_B,
                Adder64_23_in_A,
                Adder64_23_in_B,
                Adder64_24_in_A,
                Adder64_24_in_B,
                Adder64_25_in_A,
                Adder64_25_in_B,
                Adder64_26_in_A,
                Adder64_26_in_B,
                Adder64_27_in_A,
                Adder64_27_in_B,
                Adder64_28_in_A,
                Adder64_28_in_B,
                Adder64_29_in_A,
                Adder64_29_in_B,
                Adder64_30_in_A,
                Adder64_30_in_B,
                Adder64_31_in_A,
                Adder64_31_in_B,
                Adder64_32_in_A,
                Adder64_32_in_B,
                Adder64_33_in_A,
                Adder64_33_in_B,
                Adder64_34_in_A,
                Adder64_34_in_B,
                Adder64_35_in_A,
                Adder64_35_in_B,
                Adder64_36_in_A,
                Adder64_36_in_B,
                Adder64_37_in_A,
                Adder64_37_in_B,
                Adder64_38_in_A,
                Adder64_38_in_B,
                Adder64_39_in_A,
                Adder64_39_in_B,
                Adder64_40_in_A,
                Adder64_40_in_B,
                Adder64_41_in_A,
                Adder64_41_in_B,
                Adder64_42_in_A,
                Adder64_42_in_B,
                Adder64_43_in_A,
                Adder64_43_in_B,
                Adder64_44_in_A,
                Adder64_44_in_B,
                Adder64_45_in_A,
                Adder64_45_in_B,
                Adder64_46_in_A,
                Adder64_46_in_B,
                Adder64_47_in_A,
                Adder64_47_in_B,
                Adder64_48_in_A,
                Adder64_48_in_B,
                Adder64_49_in_A,
                Adder64_49_in_B,
                Adder64_50_in_A,
                Adder64_50_in_B,
                Adder64_51_in_A,
                Adder64_51_in_B,
                Adder64_52_in_A,
                Adder64_52_in_B,
                Adder64_53_in_A,
                Adder64_53_in_B,
                Adder64_54_in_A,
                Adder64_54_in_B,
                Adder64_55_in_A,
                Adder64_55_in_B,
                Adder64_56_in_A,
                Adder64_56_in_B,
                Adder64_57_in_A,
                Adder64_57_in_B,
                Adder64_58_in_A,
                Adder64_58_in_B,
                Adder64_59_in_A,
                Adder64_59_in_B,
                Adder64_60_in_A,
                Adder64_60_in_B,
                Adder64_61_in_A,
                Adder64_61_in_B,
                Adder64_62_in_A,
                Adder64_62_in_B,
                Adder64_63_in_A,
                Adder64_63_in_B,
                Adder32_0_in_A,
                Adder32_0_in_B,
                Adder32_1_in_A,
                Adder32_1_in_B,
                Adder32_2_in_A,
                Adder32_2_in_B,
                Adder32_3_in_A,
                Adder32_3_in_B,
                Adder32_4_in_A,
                Adder32_4_in_B,
                Adder32_5_in_A,
                Adder32_5_in_B,
                Adder32_6_in_A,
                Adder32_6_in_B,
                Adder32_7_in_A,
                Adder32_7_in_B,
                Adder32_8_in_A,
                Adder32_8_in_B,
                Adder32_9_in_A,
                Adder32_9_in_B,
                Adder32_10_in_A,
                Adder32_10_in_B,
                Adder32_11_in_A,
                Adder32_11_in_B,
                Adder32_12_in_A,
                Adder32_12_in_B,
                Adder32_13_in_A,
                Adder32_13_in_B,
                Adder32_14_in_A,
                Adder32_14_in_B,
                Adder32_15_in_A,
                Adder32_15_in_B,
                Adder32_16_in_A,
                Adder32_16_in_B,
                Adder32_17_in_A,
                Adder32_17_in_B,
                Adder32_18_in_A,
                Adder32_18_in_B,
                Adder32_19_in_A,
                Adder32_19_in_B,
                Adder32_20_in_A,
                Adder32_20_in_B,
                Adder32_21_in_A,
                Adder32_21_in_B,
                Adder32_22_in_A,
                Adder32_22_in_B,
                Adder32_23_in_A,
                Adder32_23_in_B,
                Adder32_24_in_A,
                Adder32_24_in_B,
                Adder32_25_in_A,
                Adder32_25_in_B,
                Adder32_26_in_A,
                Adder32_26_in_B,
                Adder32_27_in_A,
                Adder32_27_in_B,
                Adder32_28_in_A,
                Adder32_28_in_B,
                Adder32_29_in_A,
                Adder32_29_in_B,
                Adder32_30_in_A,
                Adder32_30_in_B,
                Adder32_31_in_A,
                Adder32_31_in_B,
                Adder16_0_in_A,
                Adder16_0_in_B,
                Adder16_1_in_A,
                Adder16_1_in_B,
                Adder16_2_in_A,
                Adder16_2_in_B,
                Adder16_3_in_A,
                Adder16_3_in_B,
                Adder16_4_in_A,
                Adder16_4_in_B,
                Adder16_5_in_A,
                Adder16_5_in_B,
                Adder16_6_in_A,
                Adder16_6_in_B,
                Adder16_7_in_A,
                Adder16_7_in_B,
                Adder16_8_in_A,
                Adder16_8_in_B,
                Adder16_9_in_A,
                Adder16_9_in_B,
                Adder16_10_in_A,
                Adder16_10_in_B,
                Adder16_11_in_A,
                Adder16_11_in_B,
                Adder16_12_in_A,
                Adder16_12_in_B,
                Adder16_13_in_A,
                Adder16_13_in_B,
                Adder16_14_in_A,
                Adder16_14_in_B,
                Adder16_15_in_A,
                Adder16_15_in_B,
                Adder8_0_in_A,
                Adder8_0_in_B,
                Adder8_1_in_A,
                Adder8_1_in_B,
                Adder8_2_in_A,
                Adder8_2_in_B,
                Adder8_3_in_A,
                Adder8_3_in_B,
                Adder8_4_in_A,
                Adder8_4_in_B,
                Adder8_5_in_A,
                Adder8_5_in_B,
                Adder8_6_in_A,
                Adder8_6_in_B,
                Adder8_7_in_A,
                Adder8_7_in_B,
                Adder4_0_in_A,
                Adder4_0_in_B,
                Adder4_1_in_A,
                Adder4_1_in_B,
                Adder4_2_in_A,
                Adder4_2_in_B,
                Adder4_3_in_A,
                Adder4_3_in_B,
                Adder2_0_in_A,
                Adder2_0_in_B,
                Adder2_1_in_A,
                Adder2_1_in_B,
                Adder1_0_in_A,
                Adder1_0_in_B;
    
               MassReadDataMemory MRDM_0(MemAddress, WriteData, Clk, MemWrite, MemRead, AD0_in_A, AD1_in_A, AD2_in_A, AD3_in_A, AD4_in_A, AD5_in_A, AD6_in_A, AD7_in_A, AD8_in_A, AD9_in_A, AD10_in_A, AD11_in_A, AD12_in_A, AD13_in_A, AD14_in_A, AD15_in_A, AD16_in_A, AD17_in_A, AD18_in_A, AD19_in_A, AD20_in_A, AD21_in_A, AD22_in_A, AD23_in_A, AD24_in_A, AD25_in_A, AD26_in_A, AD27_in_A, AD28_in_A, AD29_in_A, AD30_in_A, AD31_in_A, AD32_in_A, AD33_in_A, AD34_in_A, AD35_in_A, AD36_in_A, AD37_in_A, AD38_in_A, AD39_in_A, AD40_in_A, AD41_in_A, AD42_in_A, AD43_in_A, AD44_in_A, AD45_in_A, AD46_in_A, AD47_in_A, AD48_in_A, AD49_in_A, AD50_in_A, AD51_in_A, AD52_in_A, AD53_in_A, AD54_in_A, AD55_in_A, AD56_in_A, AD57_in_A, AD58_in_A, AD59_in_A, AD60_in_A, AD61_in_A, AD62_in_A, AD63_in_A, AD64_in_A, AD65_in_A, AD66_in_A, AD67_in_A, AD68_in_A, AD69_in_A, AD70_in_A, AD71_in_A, AD72_in_A, AD73_in_A, AD74_in_A, AD75_in_A, AD76_in_A, AD77_in_A, AD78_in_A, AD79_in_A, AD80_in_A, AD81_in_A, AD82_in_A, AD83_in_A, AD84_in_A, AD85_in_A, AD86_in_A, AD87_in_A, AD88_in_A, AD89_in_A, AD90_in_A, AD91_in_A, AD92_in_A, AD93_in_A, AD94_in_A, AD95_in_A, AD96_in_A, AD97_in_A, AD98_in_A, AD99_in_A, AD100_in_A, AD101_in_A, AD102_in_A, AD103_in_A, AD104_in_A, AD105_in_A, AD106_in_A, AD107_in_A, AD108_in_A, AD109_in_A, AD110_in_A, AD111_in_A, AD112_in_A, AD113_in_A, AD114_in_A, AD115_in_A, AD116_in_A, AD117_in_A, AD118_in_A, AD119_in_A, AD120_in_A, AD121_in_A, AD122_in_A, AD123_in_A, AD124_in_A, AD125_in_A, AD126_in_A, AD127_in_A, AD128_in_A, AD129_in_A, AD130_in_A, AD131_in_A, AD132_in_A, AD133_in_A, AD134_in_A, AD135_in_A, AD136_in_A, AD137_in_A, AD138_in_A, AD139_in_A, AD140_in_A, AD141_in_A, AD142_in_A, AD143_in_A, AD144_in_A, AD145_in_A, AD146_in_A, AD147_in_A, AD148_in_A, AD149_in_A, AD150_in_A, AD151_in_A, AD152_in_A, AD153_in_A, AD154_in_A, AD155_in_A, AD156_in_A, AD157_in_A, AD158_in_A, AD159_in_A, AD160_in_A, AD161_in_A, AD162_in_A, AD163_in_A, AD164_in_A, AD165_in_A, AD166_in_A, AD167_in_A, AD168_in_A, AD169_in_A, AD170_in_A, AD171_in_A, AD172_in_A, AD173_in_A, AD174_in_A, AD175_in_A, AD176_in_A, AD177_in_A, AD178_in_A, AD179_in_A, AD180_in_A, AD181_in_A, AD182_in_A, AD183_in_A, AD184_in_A, AD185_in_A, AD186_in_A, AD187_in_A, AD188_in_A, AD189_in_A, AD190_in_A, AD191_in_A, AD192_in_A, AD193_in_A, AD194_in_A, AD195_in_A, AD196_in_A, AD197_in_A, AD198_in_A, AD199_in_A, AD200_in_A, AD201_in_A, AD202_in_A, AD203_in_A, AD204_in_A, AD205_in_A, AD206_in_A, AD207_in_A, AD208_in_A, AD209_in_A, AD210_in_A, AD211_in_A, AD212_in_A, AD213_in_A, AD214_in_A, AD215_in_A, AD216_in_A, AD217_in_A, AD218_in_A, AD219_in_A, AD220_in_A, AD221_in_A, AD222_in_A, AD223_in_A, AD224_in_A, AD225_in_A, AD226_in_A, AD227_in_A, AD228_in_A, AD229_in_A, AD230_in_A, AD231_in_A, AD232_in_A, AD233_in_A, AD234_in_A, AD235_in_A, AD236_in_A, AD237_in_A, AD238_in_A, AD239_in_A, AD240_in_A, AD241_in_A, AD242_in_A, AD243_in_A, AD244_in_A, AD245_in_A, AD246_in_A, AD247_in_A, AD248_in_A, AD249_in_A, AD250_in_A, AD251_in_A, AD252_in_A, AD253_in_A, AD254_in_A, AD255_in_A);
               MassReadWindowMemory MRWM_0(WindowAddress, WriteData, Clk, MemWrite, MemRead, AD0_in_B, AD1_in_B, AD2_in_B, AD3_in_B, AD4_in_B, AD5_in_B, AD6_in_B, AD7_in_B, AD8_in_B, AD9_in_B, AD10_in_B, AD11_in_B, AD12_in_B, AD13_in_B, AD14_in_B, AD15_in_B, AD16_in_B, AD17_in_B, AD18_in_B, AD19_in_B, AD20_in_B, AD21_in_B, AD22_in_B, AD23_in_B, AD24_in_B, AD25_in_B, AD26_in_B, AD27_in_B, AD28_in_B, AD29_in_B, AD30_in_B, AD31_in_B, AD32_in_B, AD33_in_B, AD34_in_B, AD35_in_B, AD36_in_B, AD37_in_B, AD38_in_B, AD39_in_B, AD40_in_B, AD41_in_B, AD42_in_B, AD43_in_B, AD44_in_B, AD45_in_B, AD46_in_B, AD47_in_B, AD48_in_B, AD49_in_B, AD50_in_B, AD51_in_B, AD52_in_B, AD53_in_B, AD54_in_B, AD55_in_B, AD56_in_B, AD57_in_B, AD58_in_B, AD59_in_B, AD60_in_B, AD61_in_B, AD62_in_B, AD63_in_B, AD64_in_B, AD65_in_B, AD66_in_B, AD67_in_B, AD68_in_B, AD69_in_B, AD70_in_B, AD71_in_B, AD72_in_B, AD73_in_B, AD74_in_B, AD75_in_B, AD76_in_B, AD77_in_B, AD78_in_B, AD79_in_B, AD80_in_B, AD81_in_B, AD82_in_B, AD83_in_B, AD84_in_B, AD85_in_B, AD86_in_B, AD87_in_B, AD88_in_B, AD89_in_B, AD90_in_B, AD91_in_B, AD92_in_B, AD93_in_B, AD94_in_B, AD95_in_B, AD96_in_B, AD97_in_B, AD98_in_B, AD99_in_B, AD100_in_B, AD101_in_B, AD102_in_B, AD103_in_B, AD104_in_B, AD105_in_B, AD106_in_B, AD107_in_B, AD108_in_B, AD109_in_B, AD110_in_B, AD111_in_B, AD112_in_B, AD113_in_B, AD114_in_B, AD115_in_B, AD116_in_B, AD117_in_B, AD118_in_B, AD119_in_B, AD120_in_B, AD121_in_B, AD122_in_B, AD123_in_B, AD124_in_B, AD125_in_B, AD126_in_B, AD127_in_B, AD128_in_B, AD129_in_B, AD130_in_B, AD131_in_B, AD132_in_B, AD133_in_B, AD134_in_B, AD135_in_B, AD136_in_B, AD137_in_B, AD138_in_B, AD139_in_B, AD140_in_B, AD141_in_B, AD142_in_B, AD143_in_B, AD144_in_B, AD145_in_B, AD146_in_B, AD147_in_B, AD148_in_B, AD149_in_B, AD150_in_B, AD151_in_B, AD152_in_B, AD153_in_B, AD154_in_B, AD155_in_B, AD156_in_B, AD157_in_B, AD158_in_B, AD159_in_B, AD160_in_B, AD161_in_B, AD162_in_B, AD163_in_B, AD164_in_B, AD165_in_B, AD166_in_B, AD167_in_B, AD168_in_B, AD169_in_B, AD170_in_B, AD171_in_B, AD172_in_B, AD173_in_B, AD174_in_B, AD175_in_B, AD176_in_B, AD177_in_B, AD178_in_B, AD179_in_B, AD180_in_B, AD181_in_B, AD182_in_B, AD183_in_B, AD184_in_B, AD185_in_B, AD186_in_B, AD187_in_B, AD188_in_B, AD189_in_B, AD190_in_B, AD191_in_B, AD192_in_B, AD193_in_B, AD194_in_B, AD195_in_B, AD196_in_B, AD197_in_B, AD198_in_B, AD199_in_B, AD200_in_B, AD201_in_B, AD202_in_B, AD203_in_B, AD204_in_B, AD205_in_B, AD206_in_B, AD207_in_B, AD208_in_B, AD209_in_B, AD210_in_B, AD211_in_B, AD212_in_B, AD213_in_B, AD214_in_B, AD215_in_B, AD216_in_B, AD217_in_B, AD218_in_B, AD219_in_B, AD220_in_B, AD221_in_B, AD222_in_B, AD223_in_B, AD224_in_B, AD225_in_B, AD226_in_B, AD227_in_B, AD228_in_B, AD229_in_B, AD230_in_B, AD231_in_B, AD232_in_B, AD233_in_B, AD234_in_B, AD235_in_B, AD236_in_B, AD237_in_B, AD238_in_B, AD239_in_B, AD240_in_B, AD241_in_B, AD242_in_B, AD243_in_B, AD244_in_B, AD245_in_B, AD246_in_B, AD247_in_B, AD248_in_B, AD249_in_B, AD250_in_B, AD251_in_B, AD252_in_B, AD253_in_B, AD254_in_B, AD255_in_B);
                
    
                AbsoluteDifference AD0(AD0_in_A, AD0_in_B, Adder128_0_in_A);
                AbsoluteDifference AD1(AD1_in_A, AD1_in_B, Adder128_0_in_B);
                AbsoluteDifference AD2(AD2_in_A, AD2_in_B, Adder128_1_in_A);
                AbsoluteDifference AD3(AD3_in_A, AD3_in_B, Adder128_1_in_B);
                AbsoluteDifference AD4(AD4_in_A, AD4_in_B, Adder128_2_in_A);
                AbsoluteDifference AD5(AD5_in_A, AD5_in_B, Adder128_2_in_B);
                AbsoluteDifference AD6(AD6_in_A, AD6_in_B, Adder128_3_in_A);
                AbsoluteDifference AD7(AD7_in_A, AD7_in_B, Adder128_3_in_B);
                AbsoluteDifference AD8(AD8_in_A, AD8_in_B, Adder128_4_in_A);
                AbsoluteDifference AD9(AD9_in_A, AD9_in_B, Adder128_4_in_B);
                AbsoluteDifference AD10(AD10_in_A, AD10_in_B, Adder128_5_in_A);
                AbsoluteDifference AD11(AD11_in_A, AD11_in_B, Adder128_5_in_B);
                AbsoluteDifference AD12(AD12_in_A, AD12_in_B, Adder128_6_in_A);
                AbsoluteDifference AD13(AD13_in_A, AD13_in_B, Adder128_6_in_B);
                AbsoluteDifference AD14(AD14_in_A, AD14_in_B, Adder128_7_in_A);
                AbsoluteDifference AD15(AD15_in_A, AD15_in_B, Adder128_7_in_B);
                AbsoluteDifference AD16(AD16_in_A, AD16_in_B, Adder128_8_in_A);
                AbsoluteDifference AD17(AD17_in_A, AD17_in_B, Adder128_8_in_B);
                AbsoluteDifference AD18(AD18_in_A, AD18_in_B, Adder128_9_in_A);
                AbsoluteDifference AD19(AD19_in_A, AD19_in_B, Adder128_9_in_B);
                AbsoluteDifference AD20(AD20_in_A, AD20_in_B, Adder128_10_in_A);
                AbsoluteDifference AD21(AD21_in_A, AD21_in_B, Adder128_10_in_B);
                AbsoluteDifference AD22(AD22_in_A, AD22_in_B, Adder128_11_in_A);
                AbsoluteDifference AD23(AD23_in_A, AD23_in_B, Adder128_11_in_B);
                AbsoluteDifference AD24(AD24_in_A, AD24_in_B, Adder128_12_in_A);
                AbsoluteDifference AD25(AD25_in_A, AD25_in_B, Adder128_12_in_B);
                AbsoluteDifference AD26(AD26_in_A, AD26_in_B, Adder128_13_in_A);
                AbsoluteDifference AD27(AD27_in_A, AD27_in_B, Adder128_13_in_B);
                AbsoluteDifference AD28(AD28_in_A, AD28_in_B, Adder128_14_in_A);
                AbsoluteDifference AD29(AD29_in_A, AD29_in_B, Adder128_14_in_B);
                AbsoluteDifference AD30(AD30_in_A, AD30_in_B, Adder128_15_in_A);
                AbsoluteDifference AD31(AD31_in_A, AD31_in_B, Adder128_15_in_B);
                AbsoluteDifference AD32(AD32_in_A, AD32_in_B, Adder128_16_in_A);
                AbsoluteDifference AD33(AD33_in_A, AD33_in_B, Adder128_16_in_B);
                AbsoluteDifference AD34(AD34_in_A, AD34_in_B, Adder128_17_in_A);
                AbsoluteDifference AD35(AD35_in_A, AD35_in_B, Adder128_17_in_B);
                AbsoluteDifference AD36(AD36_in_A, AD36_in_B, Adder128_18_in_A);
                AbsoluteDifference AD37(AD37_in_A, AD37_in_B, Adder128_18_in_B);
                AbsoluteDifference AD38(AD38_in_A, AD38_in_B, Adder128_19_in_A);
                AbsoluteDifference AD39(AD39_in_A, AD39_in_B, Adder128_19_in_B);
                AbsoluteDifference AD40(AD40_in_A, AD40_in_B, Adder128_20_in_A);
                AbsoluteDifference AD41(AD41_in_A, AD41_in_B, Adder128_20_in_B);
                AbsoluteDifference AD42(AD42_in_A, AD42_in_B, Adder128_21_in_A);
                AbsoluteDifference AD43(AD43_in_A, AD43_in_B, Adder128_21_in_B);
                AbsoluteDifference AD44(AD44_in_A, AD44_in_B, Adder128_22_in_A);
                AbsoluteDifference AD45(AD45_in_A, AD45_in_B, Adder128_22_in_B);
                AbsoluteDifference AD46(AD46_in_A, AD46_in_B, Adder128_23_in_A);
                AbsoluteDifference AD47(AD47_in_A, AD47_in_B, Adder128_23_in_B);
                AbsoluteDifference AD48(AD48_in_A, AD48_in_B, Adder128_24_in_A);
                AbsoluteDifference AD49(AD49_in_A, AD49_in_B, Adder128_24_in_B);
                AbsoluteDifference AD50(AD50_in_A, AD50_in_B, Adder128_25_in_A);
                AbsoluteDifference AD51(AD51_in_A, AD51_in_B, Adder128_25_in_B);
                AbsoluteDifference AD52(AD52_in_A, AD52_in_B, Adder128_26_in_A);
                AbsoluteDifference AD53(AD53_in_A, AD53_in_B, Adder128_26_in_B);
                AbsoluteDifference AD54(AD54_in_A, AD54_in_B, Adder128_27_in_A);
                AbsoluteDifference AD55(AD55_in_A, AD55_in_B, Adder128_27_in_B);
                AbsoluteDifference AD56(AD56_in_A, AD56_in_B, Adder128_28_in_A);
                AbsoluteDifference AD57(AD57_in_A, AD57_in_B, Adder128_28_in_B);
                AbsoluteDifference AD58(AD58_in_A, AD58_in_B, Adder128_29_in_A);
                AbsoluteDifference AD59(AD59_in_A, AD59_in_B, Adder128_29_in_B);
                AbsoluteDifference AD60(AD60_in_A, AD60_in_B, Adder128_30_in_A);
                AbsoluteDifference AD61(AD61_in_A, AD61_in_B, Adder128_30_in_B);
                AbsoluteDifference AD62(AD62_in_A, AD62_in_B, Adder128_31_in_A);
                AbsoluteDifference AD63(AD63_in_A, AD63_in_B, Adder128_31_in_B);
                AbsoluteDifference AD64(AD64_in_A, AD64_in_B, Adder128_32_in_A);
                AbsoluteDifference AD65(AD65_in_A, AD65_in_B, Adder128_32_in_B);
                AbsoluteDifference AD66(AD66_in_A, AD66_in_B, Adder128_33_in_A);
                AbsoluteDifference AD67(AD67_in_A, AD67_in_B, Adder128_33_in_B);
                AbsoluteDifference AD68(AD68_in_A, AD68_in_B, Adder128_34_in_A);
                AbsoluteDifference AD69(AD69_in_A, AD69_in_B, Adder128_34_in_B);
                AbsoluteDifference AD70(AD70_in_A, AD70_in_B, Adder128_35_in_A);
                AbsoluteDifference AD71(AD71_in_A, AD71_in_B, Adder128_35_in_B);
                AbsoluteDifference AD72(AD72_in_A, AD72_in_B, Adder128_36_in_A);
                AbsoluteDifference AD73(AD73_in_A, AD73_in_B, Adder128_36_in_B);
                AbsoluteDifference AD74(AD74_in_A, AD74_in_B, Adder128_37_in_A);
                AbsoluteDifference AD75(AD75_in_A, AD75_in_B, Adder128_37_in_B);
                AbsoluteDifference AD76(AD76_in_A, AD76_in_B, Adder128_38_in_A);
                AbsoluteDifference AD77(AD77_in_A, AD77_in_B, Adder128_38_in_B);
                AbsoluteDifference AD78(AD78_in_A, AD78_in_B, Adder128_39_in_A);
                AbsoluteDifference AD79(AD79_in_A, AD79_in_B, Adder128_39_in_B);
                AbsoluteDifference AD80(AD80_in_A, AD80_in_B, Adder128_40_in_A);
                AbsoluteDifference AD81(AD81_in_A, AD81_in_B, Adder128_40_in_B);
                AbsoluteDifference AD82(AD82_in_A, AD82_in_B, Adder128_41_in_A);
                AbsoluteDifference AD83(AD83_in_A, AD83_in_B, Adder128_41_in_B);
                AbsoluteDifference AD84(AD84_in_A, AD84_in_B, Adder128_42_in_A);
                AbsoluteDifference AD85(AD85_in_A, AD85_in_B, Adder128_42_in_B);
                AbsoluteDifference AD86(AD86_in_A, AD86_in_B, Adder128_43_in_A);
                AbsoluteDifference AD87(AD87_in_A, AD87_in_B, Adder128_43_in_B);
                AbsoluteDifference AD88(AD88_in_A, AD88_in_B, Adder128_44_in_A);
                AbsoluteDifference AD89(AD89_in_A, AD89_in_B, Adder128_44_in_B);
                AbsoluteDifference AD90(AD90_in_A, AD90_in_B, Adder128_45_in_A);
                AbsoluteDifference AD91(AD91_in_A, AD91_in_B, Adder128_45_in_B);
                AbsoluteDifference AD92(AD92_in_A, AD92_in_B, Adder128_46_in_A);
                AbsoluteDifference AD93(AD93_in_A, AD93_in_B, Adder128_46_in_B);
                AbsoluteDifference AD94(AD94_in_A, AD94_in_B, Adder128_47_in_A);
                AbsoluteDifference AD95(AD95_in_A, AD95_in_B, Adder128_47_in_B);
                AbsoluteDifference AD96(AD96_in_A, AD96_in_B, Adder128_48_in_A);
                AbsoluteDifference AD97(AD97_in_A, AD97_in_B, Adder128_48_in_B);
                AbsoluteDifference AD98(AD98_in_A, AD98_in_B, Adder128_49_in_A);
                AbsoluteDifference AD99(AD99_in_A, AD99_in_B, Adder128_49_in_B);
                AbsoluteDifference AD100(AD100_in_A, AD100_in_B, Adder128_50_in_A);
                AbsoluteDifference AD101(AD101_in_A, AD101_in_B, Adder128_50_in_B);
                AbsoluteDifference AD102(AD102_in_A, AD102_in_B, Adder128_51_in_A);
                AbsoluteDifference AD103(AD103_in_A, AD103_in_B, Adder128_51_in_B);
                AbsoluteDifference AD104(AD104_in_A, AD104_in_B, Adder128_52_in_A);
                AbsoluteDifference AD105(AD105_in_A, AD105_in_B, Adder128_52_in_B);
                AbsoluteDifference AD106(AD106_in_A, AD106_in_B, Adder128_53_in_A);
                AbsoluteDifference AD107(AD107_in_A, AD107_in_B, Adder128_53_in_B);
                AbsoluteDifference AD108(AD108_in_A, AD108_in_B, Adder128_54_in_A);
                AbsoluteDifference AD109(AD109_in_A, AD109_in_B, Adder128_54_in_B);
                AbsoluteDifference AD110(AD110_in_A, AD110_in_B, Adder128_55_in_A);
                AbsoluteDifference AD111(AD111_in_A, AD111_in_B, Adder128_55_in_B);
                AbsoluteDifference AD112(AD112_in_A, AD112_in_B, Adder128_56_in_A);
                AbsoluteDifference AD113(AD113_in_A, AD113_in_B, Adder128_56_in_B);
                AbsoluteDifference AD114(AD114_in_A, AD114_in_B, Adder128_57_in_A);
                AbsoluteDifference AD115(AD115_in_A, AD115_in_B, Adder128_57_in_B);
                AbsoluteDifference AD116(AD116_in_A, AD116_in_B, Adder128_58_in_A);
                AbsoluteDifference AD117(AD117_in_A, AD117_in_B, Adder128_58_in_B);
                AbsoluteDifference AD118(AD118_in_A, AD118_in_B, Adder128_59_in_A);
                AbsoluteDifference AD119(AD119_in_A, AD119_in_B, Adder128_59_in_B);
                AbsoluteDifference AD120(AD120_in_A, AD120_in_B, Adder128_60_in_A);
                AbsoluteDifference AD121(AD121_in_A, AD121_in_B, Adder128_60_in_B);
                AbsoluteDifference AD122(AD122_in_A, AD122_in_B, Adder128_61_in_A);
                AbsoluteDifference AD123(AD123_in_A, AD123_in_B, Adder128_61_in_B);
                AbsoluteDifference AD124(AD124_in_A, AD124_in_B, Adder128_62_in_A);
                AbsoluteDifference AD125(AD125_in_A, AD125_in_B, Adder128_62_in_B);
                AbsoluteDifference AD126(AD126_in_A, AD126_in_B, Adder128_63_in_A);
                AbsoluteDifference AD127(AD127_in_A, AD127_in_B, Adder128_63_in_B);
                AbsoluteDifference AD128(AD128_in_A, AD128_in_B, Adder128_64_in_A);
                AbsoluteDifference AD129(AD129_in_A, AD129_in_B, Adder128_64_in_B);
                AbsoluteDifference AD130(AD130_in_A, AD130_in_B, Adder128_65_in_A);
                AbsoluteDifference AD131(AD131_in_A, AD131_in_B, Adder128_65_in_B);
                AbsoluteDifference AD132(AD132_in_A, AD132_in_B, Adder128_66_in_A);
                AbsoluteDifference AD133(AD133_in_A, AD133_in_B, Adder128_66_in_B);
                AbsoluteDifference AD134(AD134_in_A, AD134_in_B, Adder128_67_in_A);
                AbsoluteDifference AD135(AD135_in_A, AD135_in_B, Adder128_67_in_B);
                AbsoluteDifference AD136(AD136_in_A, AD136_in_B, Adder128_68_in_A);
                AbsoluteDifference AD137(AD137_in_A, AD137_in_B, Adder128_68_in_B);
                AbsoluteDifference AD138(AD138_in_A, AD138_in_B, Adder128_69_in_A);
                AbsoluteDifference AD139(AD139_in_A, AD139_in_B, Adder128_69_in_B);
                AbsoluteDifference AD140(AD140_in_A, AD140_in_B, Adder128_70_in_A);
                AbsoluteDifference AD141(AD141_in_A, AD141_in_B, Adder128_70_in_B);
                AbsoluteDifference AD142(AD142_in_A, AD142_in_B, Adder128_71_in_A);
                AbsoluteDifference AD143(AD143_in_A, AD143_in_B, Adder128_71_in_B);
                AbsoluteDifference AD144(AD144_in_A, AD144_in_B, Adder128_72_in_A);
                AbsoluteDifference AD145(AD145_in_A, AD145_in_B, Adder128_72_in_B);
                AbsoluteDifference AD146(AD146_in_A, AD146_in_B, Adder128_73_in_A);
                AbsoluteDifference AD147(AD147_in_A, AD147_in_B, Adder128_73_in_B);
                AbsoluteDifference AD148(AD148_in_A, AD148_in_B, Adder128_74_in_A);
                AbsoluteDifference AD149(AD149_in_A, AD149_in_B, Adder128_74_in_B);
                AbsoluteDifference AD150(AD150_in_A, AD150_in_B, Adder128_75_in_A);
                AbsoluteDifference AD151(AD151_in_A, AD151_in_B, Adder128_75_in_B);
                AbsoluteDifference AD152(AD152_in_A, AD152_in_B, Adder128_76_in_A);
                AbsoluteDifference AD153(AD153_in_A, AD153_in_B, Adder128_76_in_B);
                AbsoluteDifference AD154(AD154_in_A, AD154_in_B, Adder128_77_in_A);
                AbsoluteDifference AD155(AD155_in_A, AD155_in_B, Adder128_77_in_B);
                AbsoluteDifference AD156(AD156_in_A, AD156_in_B, Adder128_78_in_A);
                AbsoluteDifference AD157(AD157_in_A, AD157_in_B, Adder128_78_in_B);
                AbsoluteDifference AD158(AD158_in_A, AD158_in_B, Adder128_79_in_A);
                AbsoluteDifference AD159(AD159_in_A, AD159_in_B, Adder128_79_in_B);
                AbsoluteDifference AD160(AD160_in_A, AD160_in_B, Adder128_80_in_A);
                AbsoluteDifference AD161(AD161_in_A, AD161_in_B, Adder128_80_in_B);
                AbsoluteDifference AD162(AD162_in_A, AD162_in_B, Adder128_81_in_A);
                AbsoluteDifference AD163(AD163_in_A, AD163_in_B, Adder128_81_in_B);
                AbsoluteDifference AD164(AD164_in_A, AD164_in_B, Adder128_82_in_A);
                AbsoluteDifference AD165(AD165_in_A, AD165_in_B, Adder128_82_in_B);
                AbsoluteDifference AD166(AD166_in_A, AD166_in_B, Adder128_83_in_A);
                AbsoluteDifference AD167(AD167_in_A, AD167_in_B, Adder128_83_in_B);
                AbsoluteDifference AD168(AD168_in_A, AD168_in_B, Adder128_84_in_A);
                AbsoluteDifference AD169(AD169_in_A, AD169_in_B, Adder128_84_in_B);
                AbsoluteDifference AD170(AD170_in_A, AD170_in_B, Adder128_85_in_A);
                AbsoluteDifference AD171(AD171_in_A, AD171_in_B, Adder128_85_in_B);
                AbsoluteDifference AD172(AD172_in_A, AD172_in_B, Adder128_86_in_A);
                AbsoluteDifference AD173(AD173_in_A, AD173_in_B, Adder128_86_in_B);
                AbsoluteDifference AD174(AD174_in_A, AD174_in_B, Adder128_87_in_A);
                AbsoluteDifference AD175(AD175_in_A, AD175_in_B, Adder128_87_in_B);
                AbsoluteDifference AD176(AD176_in_A, AD176_in_B, Adder128_88_in_A);
                AbsoluteDifference AD177(AD177_in_A, AD177_in_B, Adder128_88_in_B);
                AbsoluteDifference AD178(AD178_in_A, AD178_in_B, Adder128_89_in_A);
                AbsoluteDifference AD179(AD179_in_A, AD179_in_B, Adder128_89_in_B);
                AbsoluteDifference AD180(AD180_in_A, AD180_in_B, Adder128_90_in_A);
                AbsoluteDifference AD181(AD181_in_A, AD181_in_B, Adder128_90_in_B);
                AbsoluteDifference AD182(AD182_in_A, AD182_in_B, Adder128_91_in_A);
                AbsoluteDifference AD183(AD183_in_A, AD183_in_B, Adder128_91_in_B);
                AbsoluteDifference AD184(AD184_in_A, AD184_in_B, Adder128_92_in_A);
                AbsoluteDifference AD185(AD185_in_A, AD185_in_B, Adder128_92_in_B);
                AbsoluteDifference AD186(AD186_in_A, AD186_in_B, Adder128_93_in_A);
                AbsoluteDifference AD187(AD187_in_A, AD187_in_B, Adder128_93_in_B);
                AbsoluteDifference AD188(AD188_in_A, AD188_in_B, Adder128_94_in_A);
                AbsoluteDifference AD189(AD189_in_A, AD189_in_B, Adder128_94_in_B);
                AbsoluteDifference AD190(AD190_in_A, AD190_in_B, Adder128_95_in_A);
                AbsoluteDifference AD191(AD191_in_A, AD191_in_B, Adder128_95_in_B);
                AbsoluteDifference AD192(AD192_in_A, AD192_in_B, Adder128_96_in_A);
                AbsoluteDifference AD193(AD193_in_A, AD193_in_B, Adder128_96_in_B);
                AbsoluteDifference AD194(AD194_in_A, AD194_in_B, Adder128_97_in_A);
                AbsoluteDifference AD195(AD195_in_A, AD195_in_B, Adder128_97_in_B);
                AbsoluteDifference AD196(AD196_in_A, AD196_in_B, Adder128_98_in_A);
                AbsoluteDifference AD197(AD197_in_A, AD197_in_B, Adder128_98_in_B);
                AbsoluteDifference AD198(AD198_in_A, AD198_in_B, Adder128_99_in_A);
                AbsoluteDifference AD199(AD199_in_A, AD199_in_B, Adder128_99_in_B);
                AbsoluteDifference AD200(AD200_in_A, AD200_in_B, Adder128_100_in_A);
                AbsoluteDifference AD201(AD201_in_A, AD201_in_B, Adder128_100_in_B);
                AbsoluteDifference AD202(AD202_in_A, AD202_in_B, Adder128_101_in_A);
                AbsoluteDifference AD203(AD203_in_A, AD203_in_B, Adder128_101_in_B);
                AbsoluteDifference AD204(AD204_in_A, AD204_in_B, Adder128_102_in_A);
                AbsoluteDifference AD205(AD205_in_A, AD205_in_B, Adder128_102_in_B);
                AbsoluteDifference AD206(AD206_in_A, AD206_in_B, Adder128_103_in_A);
                AbsoluteDifference AD207(AD207_in_A, AD207_in_B, Adder128_103_in_B);
                AbsoluteDifference AD208(AD208_in_A, AD208_in_B, Adder128_104_in_A);
                AbsoluteDifference AD209(AD209_in_A, AD209_in_B, Adder128_104_in_B);
                AbsoluteDifference AD210(AD210_in_A, AD210_in_B, Adder128_105_in_A);
                AbsoluteDifference AD211(AD211_in_A, AD211_in_B, Adder128_105_in_B);
                AbsoluteDifference AD212(AD212_in_A, AD212_in_B, Adder128_106_in_A);
                AbsoluteDifference AD213(AD213_in_A, AD213_in_B, Adder128_106_in_B);
                AbsoluteDifference AD214(AD214_in_A, AD214_in_B, Adder128_107_in_A);
                AbsoluteDifference AD215(AD215_in_A, AD215_in_B, Adder128_107_in_B);
                AbsoluteDifference AD216(AD216_in_A, AD216_in_B, Adder128_108_in_A);
                AbsoluteDifference AD217(AD217_in_A, AD217_in_B, Adder128_108_in_B);
                AbsoluteDifference AD218(AD218_in_A, AD218_in_B, Adder128_109_in_A);
                AbsoluteDifference AD219(AD219_in_A, AD219_in_B, Adder128_109_in_B);
                AbsoluteDifference AD220(AD220_in_A, AD220_in_B, Adder128_110_in_A);
                AbsoluteDifference AD221(AD221_in_A, AD221_in_B, Adder128_110_in_B);
                AbsoluteDifference AD222(AD222_in_A, AD222_in_B, Adder128_111_in_A);
                AbsoluteDifference AD223(AD223_in_A, AD223_in_B, Adder128_111_in_B);
                AbsoluteDifference AD224(AD224_in_A, AD224_in_B, Adder128_112_in_A);
                AbsoluteDifference AD225(AD225_in_A, AD225_in_B, Adder128_112_in_B);
                AbsoluteDifference AD226(AD226_in_A, AD226_in_B, Adder128_113_in_A);
                AbsoluteDifference AD227(AD227_in_A, AD227_in_B, Adder128_113_in_B);
                AbsoluteDifference AD228(AD228_in_A, AD228_in_B, Adder128_114_in_A);
                AbsoluteDifference AD229(AD229_in_A, AD229_in_B, Adder128_114_in_B);
                AbsoluteDifference AD230(AD230_in_A, AD230_in_B, Adder128_115_in_A);
                AbsoluteDifference AD231(AD231_in_A, AD231_in_B, Adder128_115_in_B);
                AbsoluteDifference AD232(AD232_in_A, AD232_in_B, Adder128_116_in_A);
                AbsoluteDifference AD233(AD233_in_A, AD233_in_B, Adder128_116_in_B);
                AbsoluteDifference AD234(AD234_in_A, AD234_in_B, Adder128_117_in_A);
                AbsoluteDifference AD235(AD235_in_A, AD235_in_B, Adder128_117_in_B);
                AbsoluteDifference AD236(AD236_in_A, AD236_in_B, Adder128_118_in_A);
                AbsoluteDifference AD237(AD237_in_A, AD237_in_B, Adder128_118_in_B);
                AbsoluteDifference AD238(AD238_in_A, AD238_in_B, Adder128_119_in_A);
                AbsoluteDifference AD239(AD239_in_A, AD239_in_B, Adder128_119_in_B);
                AbsoluteDifference AD240(AD240_in_A, AD240_in_B, Adder128_120_in_A);
                AbsoluteDifference AD241(AD241_in_A, AD241_in_B, Adder128_120_in_B);
                AbsoluteDifference AD242(AD242_in_A, AD242_in_B, Adder128_121_in_A);
                AbsoluteDifference AD243(AD243_in_A, AD243_in_B, Adder128_121_in_B);
                AbsoluteDifference AD244(AD244_in_A, AD244_in_B, Adder128_122_in_A);
                AbsoluteDifference AD245(AD245_in_A, AD245_in_B, Adder128_122_in_B);
                AbsoluteDifference AD246(AD246_in_A, AD246_in_B, Adder128_123_in_A);
                AbsoluteDifference AD247(AD247_in_A, AD247_in_B, Adder128_123_in_B);
                AbsoluteDifference AD248(AD248_in_A, AD248_in_B, Adder128_124_in_A);
                AbsoluteDifference AD249(AD249_in_A, AD249_in_B, Adder128_124_in_B);
                AbsoluteDifference AD250(AD250_in_A, AD250_in_B, Adder128_125_in_A);
                AbsoluteDifference AD251(AD251_in_A, AD251_in_B, Adder128_125_in_B);
                AbsoluteDifference AD252(AD252_in_A, AD252_in_B, Adder128_126_in_A);
                AbsoluteDifference AD253(AD253_in_A, AD253_in_B, Adder128_126_in_B);
                AbsoluteDifference AD254(AD254_in_A, AD254_in_B, Adder128_127_in_A);
                AbsoluteDifference AD255(AD255_in_A, AD255_in_B, Adder128_127_in_B);
    
    
                Adder Adder_128_0(Adder128_0_in_A, Adder128_0_in_B, Adder64_0_in_A);
                Adder Adder_128_1(Adder128_1_in_A, Adder128_1_in_B, Adder64_0_in_B);
                Adder Adder_128_2(Adder128_2_in_A, Adder128_2_in_B, Adder64_1_in_A);
                Adder Adder_128_3(Adder128_3_in_A, Adder128_3_in_B, Adder64_1_in_B);
                Adder Adder_128_4(Adder128_4_in_A, Adder128_4_in_B, Adder64_2_in_A);
                Adder Adder_128_5(Adder128_5_in_A, Adder128_5_in_B, Adder64_2_in_B);
                Adder Adder_128_6(Adder128_6_in_A, Adder128_6_in_B, Adder64_3_in_A);
                Adder Adder_128_7(Adder128_7_in_A, Adder128_7_in_B, Adder64_3_in_B);
                Adder Adder_128_8(Adder128_8_in_A, Adder128_8_in_B, Adder64_4_in_A);
                Adder Adder_128_9(Adder128_9_in_A, Adder128_9_in_B, Adder64_4_in_B);
                Adder Adder_128_10(Adder128_10_in_A, Adder128_10_in_B, Adder64_5_in_A);
                Adder Adder_128_11(Adder128_11_in_A, Adder128_11_in_B, Adder64_5_in_B);
                Adder Adder_128_12(Adder128_12_in_A, Adder128_12_in_B, Adder64_6_in_A);
                Adder Adder_128_13(Adder128_13_in_A, Adder128_13_in_B, Adder64_6_in_B);
                Adder Adder_128_14(Adder128_14_in_A, Adder128_14_in_B, Adder64_7_in_A);
                Adder Adder_128_15(Adder128_15_in_A, Adder128_15_in_B, Adder64_7_in_B);
                Adder Adder_128_16(Adder128_16_in_A, Adder128_16_in_B, Adder64_8_in_A);
                Adder Adder_128_17(Adder128_17_in_A, Adder128_17_in_B, Adder64_8_in_B);
                Adder Adder_128_18(Adder128_18_in_A, Adder128_18_in_B, Adder64_9_in_A);
                Adder Adder_128_19(Adder128_19_in_A, Adder128_19_in_B, Adder64_9_in_B);
                Adder Adder_128_20(Adder128_20_in_A, Adder128_20_in_B, Adder64_10_in_A);
                Adder Adder_128_21(Adder128_21_in_A, Adder128_21_in_B, Adder64_10_in_B);
                Adder Adder_128_22(Adder128_22_in_A, Adder128_22_in_B, Adder64_11_in_A);
                Adder Adder_128_23(Adder128_23_in_A, Adder128_23_in_B, Adder64_11_in_B);
                Adder Adder_128_24(Adder128_24_in_A, Adder128_24_in_B, Adder64_12_in_A);
                Adder Adder_128_25(Adder128_25_in_A, Adder128_25_in_B, Adder64_12_in_B);
                Adder Adder_128_26(Adder128_26_in_A, Adder128_26_in_B, Adder64_13_in_A);
                Adder Adder_128_27(Adder128_27_in_A, Adder128_27_in_B, Adder64_13_in_B);
                Adder Adder_128_28(Adder128_28_in_A, Adder128_28_in_B, Adder64_14_in_A);
                Adder Adder_128_29(Adder128_29_in_A, Adder128_29_in_B, Adder64_14_in_B);
                Adder Adder_128_30(Adder128_30_in_A, Adder128_30_in_B, Adder64_15_in_A);
                Adder Adder_128_31(Adder128_31_in_A, Adder128_31_in_B, Adder64_15_in_B);
                Adder Adder_128_32(Adder128_32_in_A, Adder128_32_in_B, Adder64_16_in_A);
                Adder Adder_128_33(Adder128_33_in_A, Adder128_33_in_B, Adder64_16_in_B);
                Adder Adder_128_34(Adder128_34_in_A, Adder128_34_in_B, Adder64_17_in_A);
                Adder Adder_128_35(Adder128_35_in_A, Adder128_35_in_B, Adder64_17_in_B);
                Adder Adder_128_36(Adder128_36_in_A, Adder128_36_in_B, Adder64_18_in_A);
                Adder Adder_128_37(Adder128_37_in_A, Adder128_37_in_B, Adder64_18_in_B);
                Adder Adder_128_38(Adder128_38_in_A, Adder128_38_in_B, Adder64_19_in_A);
                Adder Adder_128_39(Adder128_39_in_A, Adder128_39_in_B, Adder64_19_in_B);
                Adder Adder_128_40(Adder128_40_in_A, Adder128_40_in_B, Adder64_20_in_A);
                Adder Adder_128_41(Adder128_41_in_A, Adder128_41_in_B, Adder64_20_in_B);
                Adder Adder_128_42(Adder128_42_in_A, Adder128_42_in_B, Adder64_21_in_A);
                Adder Adder_128_43(Adder128_43_in_A, Adder128_43_in_B, Adder64_21_in_B);
                Adder Adder_128_44(Adder128_44_in_A, Adder128_44_in_B, Adder64_22_in_A);
                Adder Adder_128_45(Adder128_45_in_A, Adder128_45_in_B, Adder64_22_in_B);
                Adder Adder_128_46(Adder128_46_in_A, Adder128_46_in_B, Adder64_23_in_A);
                Adder Adder_128_47(Adder128_47_in_A, Adder128_47_in_B, Adder64_23_in_B);
                Adder Adder_128_48(Adder128_48_in_A, Adder128_48_in_B, Adder64_24_in_A);
                Adder Adder_128_49(Adder128_49_in_A, Adder128_49_in_B, Adder64_24_in_B);
                Adder Adder_128_50(Adder128_50_in_A, Adder128_50_in_B, Adder64_25_in_A);
                Adder Adder_128_51(Adder128_51_in_A, Adder128_51_in_B, Adder64_25_in_B);
                Adder Adder_128_52(Adder128_52_in_A, Adder128_52_in_B, Adder64_26_in_A);
                Adder Adder_128_53(Adder128_53_in_A, Adder128_53_in_B, Adder64_26_in_B);
                Adder Adder_128_54(Adder128_54_in_A, Adder128_54_in_B, Adder64_27_in_A);
                Adder Adder_128_55(Adder128_55_in_A, Adder128_55_in_B, Adder64_27_in_B);
                Adder Adder_128_56(Adder128_56_in_A, Adder128_56_in_B, Adder64_28_in_A);
                Adder Adder_128_57(Adder128_57_in_A, Adder128_57_in_B, Adder64_28_in_B);
                Adder Adder_128_58(Adder128_58_in_A, Adder128_58_in_B, Adder64_29_in_A);
                Adder Adder_128_59(Adder128_59_in_A, Adder128_59_in_B, Adder64_29_in_B);
                Adder Adder_128_60(Adder128_60_in_A, Adder128_60_in_B, Adder64_30_in_A);
                Adder Adder_128_61(Adder128_61_in_A, Adder128_61_in_B, Adder64_30_in_B);
                Adder Adder_128_62(Adder128_62_in_A, Adder128_62_in_B, Adder64_31_in_A);
                Adder Adder_128_63(Adder128_63_in_A, Adder128_63_in_B, Adder64_31_in_B);
                Adder Adder_128_64(Adder128_64_in_A, Adder128_64_in_B, Adder64_32_in_A);
                Adder Adder_128_65(Adder128_65_in_A, Adder128_65_in_B, Adder64_32_in_B);
                Adder Adder_128_66(Adder128_66_in_A, Adder128_66_in_B, Adder64_33_in_A);
                Adder Adder_128_67(Adder128_67_in_A, Adder128_67_in_B, Adder64_33_in_B);
                Adder Adder_128_68(Adder128_68_in_A, Adder128_68_in_B, Adder64_34_in_A);
                Adder Adder_128_69(Adder128_69_in_A, Adder128_69_in_B, Adder64_34_in_B);
                Adder Adder_128_70(Adder128_70_in_A, Adder128_70_in_B, Adder64_35_in_A);
                Adder Adder_128_71(Adder128_71_in_A, Adder128_71_in_B, Adder64_35_in_B);
                Adder Adder_128_72(Adder128_72_in_A, Adder128_72_in_B, Adder64_36_in_A);
                Adder Adder_128_73(Adder128_73_in_A, Adder128_73_in_B, Adder64_36_in_B);
                Adder Adder_128_74(Adder128_74_in_A, Adder128_74_in_B, Adder64_37_in_A);
                Adder Adder_128_75(Adder128_75_in_A, Adder128_75_in_B, Adder64_37_in_B);
                Adder Adder_128_76(Adder128_76_in_A, Adder128_76_in_B, Adder64_38_in_A);
                Adder Adder_128_77(Adder128_77_in_A, Adder128_77_in_B, Adder64_38_in_B);
                Adder Adder_128_78(Adder128_78_in_A, Adder128_78_in_B, Adder64_39_in_A);
                Adder Adder_128_79(Adder128_79_in_A, Adder128_79_in_B, Adder64_39_in_B);
                Adder Adder_128_80(Adder128_80_in_A, Adder128_80_in_B, Adder64_40_in_A);
                Adder Adder_128_81(Adder128_81_in_A, Adder128_81_in_B, Adder64_40_in_B);
                Adder Adder_128_82(Adder128_82_in_A, Adder128_82_in_B, Adder64_41_in_A);
                Adder Adder_128_83(Adder128_83_in_A, Adder128_83_in_B, Adder64_41_in_B);
                Adder Adder_128_84(Adder128_84_in_A, Adder128_84_in_B, Adder64_42_in_A);
                Adder Adder_128_85(Adder128_85_in_A, Adder128_85_in_B, Adder64_42_in_B);
                Adder Adder_128_86(Adder128_86_in_A, Adder128_86_in_B, Adder64_43_in_A);
                Adder Adder_128_87(Adder128_87_in_A, Adder128_87_in_B, Adder64_43_in_B);
                Adder Adder_128_88(Adder128_88_in_A, Adder128_88_in_B, Adder64_44_in_A);
                Adder Adder_128_89(Adder128_89_in_A, Adder128_89_in_B, Adder64_44_in_B);
                Adder Adder_128_90(Adder128_90_in_A, Adder128_90_in_B, Adder64_45_in_A);
                Adder Adder_128_91(Adder128_91_in_A, Adder128_91_in_B, Adder64_45_in_B);
                Adder Adder_128_92(Adder128_92_in_A, Adder128_92_in_B, Adder64_46_in_A);
                Adder Adder_128_93(Adder128_93_in_A, Adder128_93_in_B, Adder64_46_in_B);
                Adder Adder_128_94(Adder128_94_in_A, Adder128_94_in_B, Adder64_47_in_A);
                Adder Adder_128_95(Adder128_95_in_A, Adder128_95_in_B, Adder64_47_in_B);
                Adder Adder_128_96(Adder128_96_in_A, Adder128_96_in_B, Adder64_48_in_A);
                Adder Adder_128_97(Adder128_97_in_A, Adder128_97_in_B, Adder64_48_in_B);
                Adder Adder_128_98(Adder128_98_in_A, Adder128_98_in_B, Adder64_49_in_A);
                Adder Adder_128_99(Adder128_99_in_A, Adder128_99_in_B, Adder64_49_in_B);
                Adder Adder_128_100(Adder128_100_in_A, Adder128_100_in_B, Adder64_50_in_A);
                Adder Adder_128_101(Adder128_101_in_A, Adder128_101_in_B, Adder64_50_in_B);
                Adder Adder_128_102(Adder128_102_in_A, Adder128_102_in_B, Adder64_51_in_A);
                Adder Adder_128_103(Adder128_103_in_A, Adder128_103_in_B, Adder64_51_in_B);
                Adder Adder_128_104(Adder128_104_in_A, Adder128_104_in_B, Adder64_52_in_A);
                Adder Adder_128_105(Adder128_105_in_A, Adder128_105_in_B, Adder64_52_in_B);
                Adder Adder_128_106(Adder128_106_in_A, Adder128_106_in_B, Adder64_53_in_A);
                Adder Adder_128_107(Adder128_107_in_A, Adder128_107_in_B, Adder64_53_in_B);
                Adder Adder_128_108(Adder128_108_in_A, Adder128_108_in_B, Adder64_54_in_A);
                Adder Adder_128_109(Adder128_109_in_A, Adder128_109_in_B, Adder64_54_in_B);
                Adder Adder_128_110(Adder128_110_in_A, Adder128_110_in_B, Adder64_55_in_A);
                Adder Adder_128_111(Adder128_111_in_A, Adder128_111_in_B, Adder64_55_in_B);
                Adder Adder_128_112(Adder128_112_in_A, Adder128_112_in_B, Adder64_56_in_A);
                Adder Adder_128_113(Adder128_113_in_A, Adder128_113_in_B, Adder64_56_in_B);
                Adder Adder_128_114(Adder128_114_in_A, Adder128_114_in_B, Adder64_57_in_A);
                Adder Adder_128_115(Adder128_115_in_A, Adder128_115_in_B, Adder64_57_in_B);
                Adder Adder_128_116(Adder128_116_in_A, Adder128_116_in_B, Adder64_58_in_A);
                Adder Adder_128_117(Adder128_117_in_A, Adder128_117_in_B, Adder64_58_in_B);
                Adder Adder_128_118(Adder128_118_in_A, Adder128_118_in_B, Adder64_59_in_A);
                Adder Adder_128_119(Adder128_119_in_A, Adder128_119_in_B, Adder64_59_in_B);
                Adder Adder_128_120(Adder128_120_in_A, Adder128_120_in_B, Adder64_60_in_A);
                Adder Adder_128_121(Adder128_121_in_A, Adder128_121_in_B, Adder64_60_in_B);
                Adder Adder_128_122(Adder128_122_in_A, Adder128_122_in_B, Adder64_61_in_A);
                Adder Adder_128_123(Adder128_123_in_A, Adder128_123_in_B, Adder64_61_in_B);
                Adder Adder_128_124(Adder128_124_in_A, Adder128_124_in_B, Adder64_62_in_A);
                Adder Adder_128_125(Adder128_125_in_A, Adder128_125_in_B, Adder64_62_in_B);
                Adder Adder_128_126(Adder128_126_in_A, Adder128_126_in_B, Adder64_63_in_A);
                Adder Adder_128_127(Adder128_127_in_A, Adder128_127_in_B, Adder64_63_in_B);
                Adder Adder_64_0(Adder64_0_in_A, Adder64_0_in_B, Adder32_0_in_A);
                Adder Adder_64_1(Adder64_1_in_A, Adder64_1_in_B, Adder32_0_in_B);
                Adder Adder_64_2(Adder64_2_in_A, Adder64_2_in_B, Adder32_1_in_A);
                Adder Adder_64_3(Adder64_3_in_A, Adder64_3_in_B, Adder32_1_in_B);
                Adder Adder_64_4(Adder64_4_in_A, Adder64_4_in_B, Adder32_2_in_A);
                Adder Adder_64_5(Adder64_5_in_A, Adder64_5_in_B, Adder32_2_in_B);
                Adder Adder_64_6(Adder64_6_in_A, Adder64_6_in_B, Adder32_3_in_A);
                Adder Adder_64_7(Adder64_7_in_A, Adder64_7_in_B, Adder32_3_in_B);
                Adder Adder_64_8(Adder64_8_in_A, Adder64_8_in_B, Adder32_4_in_A);
                Adder Adder_64_9(Adder64_9_in_A, Adder64_9_in_B, Adder32_4_in_B);
                Adder Adder_64_10(Adder64_10_in_A, Adder64_10_in_B, Adder32_5_in_A);
                Adder Adder_64_11(Adder64_11_in_A, Adder64_11_in_B, Adder32_5_in_B);
                Adder Adder_64_12(Adder64_12_in_A, Adder64_12_in_B, Adder32_6_in_A);
                Adder Adder_64_13(Adder64_13_in_A, Adder64_13_in_B, Adder32_6_in_B);
                Adder Adder_64_14(Adder64_14_in_A, Adder64_14_in_B, Adder32_7_in_A);
                Adder Adder_64_15(Adder64_15_in_A, Adder64_15_in_B, Adder32_7_in_B);
                Adder Adder_64_16(Adder64_16_in_A, Adder64_16_in_B, Adder32_8_in_A);
                Adder Adder_64_17(Adder64_17_in_A, Adder64_17_in_B, Adder32_8_in_B);
                Adder Adder_64_18(Adder64_18_in_A, Adder64_18_in_B, Adder32_9_in_A);
                Adder Adder_64_19(Adder64_19_in_A, Adder64_19_in_B, Adder32_9_in_B);
                Adder Adder_64_20(Adder64_20_in_A, Adder64_20_in_B, Adder32_10_in_A);
                Adder Adder_64_21(Adder64_21_in_A, Adder64_21_in_B, Adder32_10_in_B);
                Adder Adder_64_22(Adder64_22_in_A, Adder64_22_in_B, Adder32_11_in_A);
                Adder Adder_64_23(Adder64_23_in_A, Adder64_23_in_B, Adder32_11_in_B);
                Adder Adder_64_24(Adder64_24_in_A, Adder64_24_in_B, Adder32_12_in_A);
                Adder Adder_64_25(Adder64_25_in_A, Adder64_25_in_B, Adder32_12_in_B);
                Adder Adder_64_26(Adder64_26_in_A, Adder64_26_in_B, Adder32_13_in_A);
                Adder Adder_64_27(Adder64_27_in_A, Adder64_27_in_B, Adder32_13_in_B);
                Adder Adder_64_28(Adder64_28_in_A, Adder64_28_in_B, Adder32_14_in_A);
                Adder Adder_64_29(Adder64_29_in_A, Adder64_29_in_B, Adder32_14_in_B);
                Adder Adder_64_30(Adder64_30_in_A, Adder64_30_in_B, Adder32_15_in_A);
                Adder Adder_64_31(Adder64_31_in_A, Adder64_31_in_B, Adder32_15_in_B);
                Adder Adder_64_32(Adder64_32_in_A, Adder64_32_in_B, Adder32_16_in_A);
                Adder Adder_64_33(Adder64_33_in_A, Adder64_33_in_B, Adder32_16_in_B);
                Adder Adder_64_34(Adder64_34_in_A, Adder64_34_in_B, Adder32_17_in_A);
                Adder Adder_64_35(Adder64_35_in_A, Adder64_35_in_B, Adder32_17_in_B);
                Adder Adder_64_36(Adder64_36_in_A, Adder64_36_in_B, Adder32_18_in_A);
                Adder Adder_64_37(Adder64_37_in_A, Adder64_37_in_B, Adder32_18_in_B);
                Adder Adder_64_38(Adder64_38_in_A, Adder64_38_in_B, Adder32_19_in_A);
                Adder Adder_64_39(Adder64_39_in_A, Adder64_39_in_B, Adder32_19_in_B);
                Adder Adder_64_40(Adder64_40_in_A, Adder64_40_in_B, Adder32_20_in_A);
                Adder Adder_64_41(Adder64_41_in_A, Adder64_41_in_B, Adder32_20_in_B);
                Adder Adder_64_42(Adder64_42_in_A, Adder64_42_in_B, Adder32_21_in_A);
                Adder Adder_64_43(Adder64_43_in_A, Adder64_43_in_B, Adder32_21_in_B);
                Adder Adder_64_44(Adder64_44_in_A, Adder64_44_in_B, Adder32_22_in_A);
                Adder Adder_64_45(Adder64_45_in_A, Adder64_45_in_B, Adder32_22_in_B);
                Adder Adder_64_46(Adder64_46_in_A, Adder64_46_in_B, Adder32_23_in_A);
                Adder Adder_64_47(Adder64_47_in_A, Adder64_47_in_B, Adder32_23_in_B);
                Adder Adder_64_48(Adder64_48_in_A, Adder64_48_in_B, Adder32_24_in_A);
                Adder Adder_64_49(Adder64_49_in_A, Adder64_49_in_B, Adder32_24_in_B);
                Adder Adder_64_50(Adder64_50_in_A, Adder64_50_in_B, Adder32_25_in_A);
                Adder Adder_64_51(Adder64_51_in_A, Adder64_51_in_B, Adder32_25_in_B);
                Adder Adder_64_52(Adder64_52_in_A, Adder64_52_in_B, Adder32_26_in_A);
                Adder Adder_64_53(Adder64_53_in_A, Adder64_53_in_B, Adder32_26_in_B);
                Adder Adder_64_54(Adder64_54_in_A, Adder64_54_in_B, Adder32_27_in_A);
                Adder Adder_64_55(Adder64_55_in_A, Adder64_55_in_B, Adder32_27_in_B);
                Adder Adder_64_56(Adder64_56_in_A, Adder64_56_in_B, Adder32_28_in_A);
                Adder Adder_64_57(Adder64_57_in_A, Adder64_57_in_B, Adder32_28_in_B);
                Adder Adder_64_58(Adder64_58_in_A, Adder64_58_in_B, Adder32_29_in_A);
                Adder Adder_64_59(Adder64_59_in_A, Adder64_59_in_B, Adder32_29_in_B);
                Adder Adder_64_60(Adder64_60_in_A, Adder64_60_in_B, Adder32_30_in_A);
                Adder Adder_64_61(Adder64_61_in_A, Adder64_61_in_B, Adder32_30_in_B);
                Adder Adder_64_62(Adder64_62_in_A, Adder64_62_in_B, Adder32_31_in_A);
                Adder Adder_64_63(Adder64_63_in_A, Adder64_63_in_B, Adder32_31_in_B);
                Adder Adder_32_0(Adder32_0_in_A, Adder32_0_in_B, Adder16_0_in_A);
                Adder Adder_32_1(Adder32_1_in_A, Adder32_1_in_B, Adder16_0_in_B);
                Adder Adder_32_2(Adder32_2_in_A, Adder32_2_in_B, Adder16_1_in_A);
                Adder Adder_32_3(Adder32_3_in_A, Adder32_3_in_B, Adder16_1_in_B);
                Adder Adder_32_4(Adder32_4_in_A, Adder32_4_in_B, Adder16_2_in_A);
                Adder Adder_32_5(Adder32_5_in_A, Adder32_5_in_B, Adder16_2_in_B);
                Adder Adder_32_6(Adder32_6_in_A, Adder32_6_in_B, Adder16_3_in_A);
                Adder Adder_32_7(Adder32_7_in_A, Adder32_7_in_B, Adder16_3_in_B);
                Adder Adder_32_8(Adder32_8_in_A, Adder32_8_in_B, Adder16_4_in_A);
                Adder Adder_32_9(Adder32_9_in_A, Adder32_9_in_B, Adder16_4_in_B);
                Adder Adder_32_10(Adder32_10_in_A, Adder32_10_in_B, Adder16_5_in_A);
                Adder Adder_32_11(Adder32_11_in_A, Adder32_11_in_B, Adder16_5_in_B);
                Adder Adder_32_12(Adder32_12_in_A, Adder32_12_in_B, Adder16_6_in_A);
                Adder Adder_32_13(Adder32_13_in_A, Adder32_13_in_B, Adder16_6_in_B);
                Adder Adder_32_14(Adder32_14_in_A, Adder32_14_in_B, Adder16_7_in_A);
                Adder Adder_32_15(Adder32_15_in_A, Adder32_15_in_B, Adder16_7_in_B);
                Adder Adder_32_16(Adder32_16_in_A, Adder32_16_in_B, Adder16_8_in_A);
                Adder Adder_32_17(Adder32_17_in_A, Adder32_17_in_B, Adder16_8_in_B);
                Adder Adder_32_18(Adder32_18_in_A, Adder32_18_in_B, Adder16_9_in_A);
                Adder Adder_32_19(Adder32_19_in_A, Adder32_19_in_B, Adder16_9_in_B);
                Adder Adder_32_20(Adder32_20_in_A, Adder32_20_in_B, Adder16_10_in_A);
                Adder Adder_32_21(Adder32_21_in_A, Adder32_21_in_B, Adder16_10_in_B);
                Adder Adder_32_22(Adder32_22_in_A, Adder32_22_in_B, Adder16_11_in_A);
                Adder Adder_32_23(Adder32_23_in_A, Adder32_23_in_B, Adder16_11_in_B);
                Adder Adder_32_24(Adder32_24_in_A, Adder32_24_in_B, Adder16_12_in_A);
                Adder Adder_32_25(Adder32_25_in_A, Adder32_25_in_B, Adder16_12_in_B);
                Adder Adder_32_26(Adder32_26_in_A, Adder32_26_in_B, Adder16_13_in_A);
                Adder Adder_32_27(Adder32_27_in_A, Adder32_27_in_B, Adder16_13_in_B);
                Adder Adder_32_28(Adder32_28_in_A, Adder32_28_in_B, Adder16_14_in_A);
                Adder Adder_32_29(Adder32_29_in_A, Adder32_29_in_B, Adder16_14_in_B);
                Adder Adder_32_30(Adder32_30_in_A, Adder32_30_in_B, Adder16_15_in_A);
                Adder Adder_32_31(Adder32_31_in_A, Adder32_31_in_B, Adder16_15_in_B);
                Adder Adder_16_0(Adder16_0_in_A, Adder16_0_in_B, Adder8_0_in_A);
                Adder Adder_16_1(Adder16_1_in_A, Adder16_1_in_B, Adder8_0_in_B);
                Adder Adder_16_2(Adder16_2_in_A, Adder16_2_in_B, Adder8_1_in_A);
                Adder Adder_16_3(Adder16_3_in_A, Adder16_3_in_B, Adder8_1_in_B);
                Adder Adder_16_4(Adder16_4_in_A, Adder16_4_in_B, Adder8_2_in_A);
                Adder Adder_16_5(Adder16_5_in_A, Adder16_5_in_B, Adder8_2_in_B);
                Adder Adder_16_6(Adder16_6_in_A, Adder16_6_in_B, Adder8_3_in_A);
                Adder Adder_16_7(Adder16_7_in_A, Adder16_7_in_B, Adder8_3_in_B);
                Adder Adder_16_8(Adder16_8_in_A, Adder16_8_in_B, Adder8_4_in_A);
                Adder Adder_16_9(Adder16_9_in_A, Adder16_9_in_B, Adder8_4_in_B);
                Adder Adder_16_10(Adder16_10_in_A, Adder16_10_in_B, Adder8_5_in_A);
                Adder Adder_16_11(Adder16_11_in_A, Adder16_11_in_B, Adder8_5_in_B);
                Adder Adder_16_12(Adder16_12_in_A, Adder16_12_in_B, Adder8_6_in_A);
                Adder Adder_16_13(Adder16_13_in_A, Adder16_13_in_B, Adder8_6_in_B);
                Adder Adder_16_14(Adder16_14_in_A, Adder16_14_in_B, Adder8_7_in_A);
                Adder Adder_16_15(Adder16_15_in_A, Adder16_15_in_B, Adder8_7_in_B);
                Adder Adder_8_0(Adder8_0_in_A, Adder8_0_in_B, Adder4_0_in_A);
                Adder Adder_8_1(Adder8_1_in_A, Adder8_1_in_B, Adder4_0_in_B);
                Adder Adder_8_2(Adder8_2_in_A, Adder8_2_in_B, Adder4_1_in_A);
                Adder Adder_8_3(Adder8_3_in_A, Adder8_3_in_B, Adder4_1_in_B);
                Adder Adder_8_4(Adder8_4_in_A, Adder8_4_in_B, Adder4_2_in_A);
                Adder Adder_8_5(Adder8_5_in_A, Adder8_5_in_B, Adder4_2_in_B);
                Adder Adder_8_6(Adder8_6_in_A, Adder8_6_in_B, Adder4_3_in_A);
                Adder Adder_8_7(Adder8_7_in_A, Adder8_7_in_B, Adder4_3_in_B);
                Adder Adder_4_0(Adder4_0_in_A, Adder4_0_in_B, Adder2_0_in_A);
                Adder Adder_4_1(Adder4_1_in_A, Adder4_1_in_B, Adder2_0_in_B);
                Adder Adder_4_2(Adder4_2_in_A, Adder4_2_in_B, Adder2_1_in_A);
                Adder Adder_4_3(Adder4_3_in_A, Adder4_3_in_B, Adder2_1_in_B);
                Adder Adder_2_0(Adder2_0_in_A, Adder2_0_in_B, Adder1_0_in_A);
                Adder Adder_2_1(Adder2_1_in_A, Adder2_1_in_B, Adder1_0_in_B);
                Adder Adder_1_0(Adder1_0_in_A, Adder1_0_in_B, SAD_out);  
    
    
endmodule
