`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/30/2018 06:01:28 PM
// Design Name: 
// Module Name: SadRegister
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SadRegister( MemWidth,  MemHeight,  FrameWidth );

    input [31:0] MemWidth, //Amount of memory per row read
                          MemHeight, //Amount of rows to read
                          FrameWidth; //width of the overall image frame

endmodule
