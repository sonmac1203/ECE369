`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369A - Computer Architecture
// Laboratory  1
// Module - InstructionMemory.v
// Description - 32-Bit wide instruction memory.
//
// INPUT:-
// Address: 32-Bit address input port.
//
// OUTPUT:-
// Instruction: 32-Bit output port.
//
// FUNCTIONALITY:-
// Similar to the DataMemory, this module should also be byte-addressed
// (i.e., ignore bits 0 and 1 of 'Address'). All of the instructions will be 
// hard-coded into the instruction memory, so there is no need to write to the 
// InstructionMemory.  The contents of the InstructionMemory is the machine 
// language program to be run on your MIPS processor.
//
//
//we will store the machine code for a code written in C later. for now initialize 
//each entry to be its index * 3 (memory[i] = i * 3;)
//all you need to do is give an address as input and read the contents of the 
//address on your output port. 
// 
//Using a 32bit address you will index into the memory, output the contents of that specific 
//address. for data memory we are using 1K word of storage space. for the instruction memory 
//you may assume smaller size for practical purpose. you can use 128 words as the size and 
//hardcode the values.  in this case you need 7 bits to index into the memory. 
//
//be careful with the least two significant bits of the 32bit address. those help us index 
//into one of the 4 bytes in a word. therefore you will need to use bit [8-2] of the input address. 


////////////////////////////////////////////////////////////////////////////////

module InstructionMemory(Address, Instruction); 

    input [31:0] Address;        // Input Address 

    output reg [31:0] Instruction;    // Instruction at memory location Address
    
    reg [31:0] memory [0:1023];

    //initializing memory with 0-127    
    //integer index;
    
    
    initial begin





memory[0] <= 32'h23bdfffc;	//	main:			addi	$sp, $sp, -4
memory[1] <= 32'hafbf0000;	//				sw	$ra, 0($sp)
memory[2] <= 32'h34040000;	//				ori	$a0, $zero, 0
memory[3] <= 32'h34050010;	//				ori	$a1, $zero, 16
memory[4] <= 32'h34060410;	//				ori	$a2, $zero, 1040
memory[5] <= 32'h0c00000a;	//				jal	vbsme
memory[6] <= 32'h0c000008;	//				jal	print_result
memory[7] <= 32'h08000007;	//	exit:			j	exit
memory[8] <= 32'h00000000;	//	print_result:		nop
memory[9] <= 32'h03e00008;	//				jr	$ra
memory[10] <= 32'h8c900000;	//	vbsme:			lw	$s0, 0($a0)
memory[11] <= 32'h8c910004;	//				lw	$s1, 4($a0)
memory[12] <= 32'h8c920008;	//				lw	$s2, 8($a0)
memory[13] <= 32'h8c93000c;	//				lw	$s3, 12($a0)
memory[14] <= 32'h340e0000;	//				ori	$t6, $zero, 0
memory[15] <= 32'h340f0000;	//				ori	$t7, $zero, 0
memory[16] <= 32'h02124022;	//				sub	$t0, $s0, $s2
memory[17] <= 32'h71114002;	//				mul	$t0, $t0, $s1
memory[18] <= 32'h02334822;	//				sub	$t1, $s1, $s3
memory[19] <= 32'h0109a820;	//				add	$s5, $t0, $t1
memory[20] <= 32'hafa80004;	//				sw	$t0, 4($sp)
memory[21] <= 32'h34020000;	//				ori	$v0, $zero, 0
memory[22] <= 32'h34030000;	//				ori	$v1, $zero, 0
memory[23] <= 32'h3416270f;	//				ori	$s6, $zero, 9999
memory[24] <= 32'h23bdfffc;	//				addi	$sp, $sp, -4
memory[25] <= 32'hafbf0000;	//				sw	$ra, 0($sp)
memory[26] <= 32'h0271402a;	//				slt	$t0, $s3, $s1
memory[27] <= 32'h0250482a;	//				slt	$t1, $s2, $s0
memory[28] <= 32'h01094025;	//				or	$t0, $t0, $t1
memory[29] <= 32'h1100003c;	//				beq	$t0, $0, endzigzag
memory[30] <= 32'h0c00005e;	//				jal	sad
memory[31] <= 32'h02334022;	//				sub	$t0, $s1, $s3
memory[32] <= 32'h01e8402a;	//				slt	$t0, $t7, $t0
memory[33] <= 32'h11000002;	//				beq	$t0, $0, errordetectnexta
memory[34] <= 32'h0c000083;	//				jal	rightsubroutine
memory[35] <= 32'h08000028;	//				j	doneerrordetectright
memory[36] <= 32'h02124022;	//	errordetectnexta:	sub	$t0, $s0, $s2
memory[37] <= 32'h01c8402a;	//				slt	$t0, $t6, $t0
memory[38] <= 32'h11000033;	//				beq	$t0, $0, endzigzag
memory[39] <= 32'h0c00008b;	//				jal	downsubroutine
memory[40] <= 32'h0c00005e;	//	doneerrordetectright:	jal	sad
memory[41] <= 32'h71d14002;	//	zigzagloop:		mul	$t0, $t6, $s1
memory[42] <= 32'h010f4020;	//				add	$t0, $t0, $t7
memory[43] <= 32'h0115402a;	//				slt	$t0, $t0, $s5
memory[44] <= 32'h1100002d;	//				beq	$t0, $0, endzigzag
memory[45] <= 32'h20140001;	//				addi	$s4, $0, 1
memory[46] <= 32'h1280000e;	//	dlcollisiondetect:	beq	$s4, $0, edlcollisiondetect
memory[47] <= 32'h02124022;	//				sub	$t0, $s0, $s2
memory[48] <= 32'h01c8402a;	//				slt	$t0, $t6, $t0
memory[49] <= 32'h11000007;	//				beq	$t0, $0, downcollisiona
memory[50] <= 32'h000f402a;	//				slt	$t0, $0, $t7
memory[51] <= 32'h11000002;	//				beq	$t0, $0, leftcollisiona
memory[52] <= 32'h0c000085;	//				jal	downleftsubroutine
memory[53] <= 32'h0800003b;	//				j	downcollisionaend
memory[54] <= 32'h0c00008b;	//	leftcollisiona:		jal	downsubroutine
memory[55] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[56] <= 32'h0800003b;	//				j	downcollisionaend
memory[57] <= 32'h0c000083;	//	downcollisiona:		jal	rightsubroutine
memory[58] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[59] <= 32'h0c00005e;	//	downcollisionaend:	jal	sad
memory[60] <= 32'h0800002e;	//				j	dlcollisiondetect
memory[61] <= 32'h0c00005e;	//	edlcollisiondetect:	jal	sad
memory[62] <= 32'h71d14002;	//				mul	$t0, $t6, $s1
memory[63] <= 32'h010f4020;	//				add	$t0, $t0, $t7
memory[64] <= 32'h0115402a;	//				slt	$t0, $t0, $s5
memory[65] <= 32'h11000018;	//				beq	$t0, $0, endzigzag
memory[66] <= 32'h20140001;	//				addi	$s4, $0, 1
memory[67] <= 32'h12800014;	//	urcollisiondetect:	beq	$s4, $0, eurcollisiondetect
memory[68] <= 32'h000e402a;	//				slt	$t0, $0, $t6
memory[69] <= 32'h11000008;	//				beq	$t0, $0, upcollisiona
memory[70] <= 32'h02334022;	//				sub	$t0, $s1, $s3
memory[71] <= 32'h01e8402a;	//				slt	$t0, $t7, $t0
memory[72] <= 32'h11000002;	//				beq	$t0, $0, rightcollisiona
memory[73] <= 32'h0c000088;	//				jal	uprightsubroutine
memory[74] <= 32'h08000056;	//				j	upcollisionaend
memory[75] <= 32'h0c00008b;	//	rightcollisiona:	jal	downsubroutine
memory[76] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[77] <= 32'h08000056;	//				j	upcollisionaend
memory[78] <= 32'h02334022;	//	upcollisiona:		sub	$t0, $s1, $s3
memory[79] <= 32'h01e8402a;	//				slt	$t0, $t7, $t0
memory[80] <= 32'h11000003;	//				beq	$t0, $0, rightcollisionb
memory[81] <= 32'h0c000083;	//				jal	rightsubroutine
memory[82] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[83] <= 32'h08000056;	//				j	upcollisionaend
memory[84] <= 32'h0c00008b;	//	rightcollisionb:	jal	downsubroutine
memory[85] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[86] <= 32'h0c00005e;	//	upcollisionaend:	jal	sad
memory[87] <= 32'h08000043;	//				j	urcollisiondetect
memory[88] <= 32'h0c00005e;	//	eurcollisiondetect:	jal	sad
memory[89] <= 32'h08000029;	//				j	zigzagloop
memory[90] <= 32'h8fbf0000;	//	endzigzag:		lw	$ra, 0($sp)
memory[91] <= 32'h00000000;	//				nop
memory[92] <= 32'h00000000;	//				nop
memory[93] <= 32'h03e00008;	//				jr	$ra
memory[94] <= 32'h00000000;	//	sad:			nop
memory[95] <= 32'h00004020;	//				add	$t0, $0, $0
memory[96] <= 32'h00004820;	//				add	$t1, $0, $0
memory[97] <= 32'h0132582a;	//	sadouterloop:		slt	$t3, $t1, $s2
memory[98] <= 32'h11600019;	//				beq	$t3, $0, sadouterloopend
memory[99] <= 32'h00005020;	//				add	$t2, $0, $0
memory[100] <= 32'h0153582a;	//	sadinnerloop:		slt	$t3, $t2, $s3
memory[101] <= 32'h11600014;	//				beq	$t3, $0, sadinnerloopend
memory[102] <= 32'h012e5820;	//				add	$t3, $t1, $t6
memory[103] <= 32'h71715802;	//				mul	$t3, $t3, $s1
memory[104] <= 32'h016a5820;	//				add	$t3, $t3, $t2
memory[105] <= 32'h016f5820;	//				add	$t3, $t3, $t7
memory[106] <= 32'h000b5880;	//				sll	$t3, $t3, 2
memory[107] <= 32'h71336002;	//				mul	$t4, $t1, $s3
memory[108] <= 32'h018a6020;	//				add	$t4, $t4, $t2
memory[109] <= 32'h000c6080;	//				sll	$t4, $t4, 2
memory[110] <= 32'h00ab5820;	//				add	$t3, $a1, $t3
memory[111] <= 32'h00cc6020;	//				add	$t4, $a2, $t4
memory[112] <= 32'h8d6b0000;	//				lw	$t3, 0($t3)
memory[113] <= 32'h8d8c0000;	//				lw	$t4, 0($t4)
memory[114] <= 32'h016c5822;	//				sub	$t3, $t3, $t4
memory[115] <= 32'h0160602a;	//				slt	$t4, $t3, $0
memory[116] <= 32'h11800002;	//				beq	$t4, $0, absifend
memory[117] <= 32'h200dffff;	//				addi	$t5, $0, -1
memory[118] <= 32'h716d5802;	//				mul	$t3, $t3, $t5
memory[119] <= 32'h010b4020;	//	absifend:		add	$t0, $t0, $t3
memory[120] <= 32'h214a0001;	//				addi	$t2, $t2, 1
memory[121] <= 32'h08000064;	//				j	sadinnerloop
memory[122] <= 32'h21290001;	//	sadinnerloopend:	addi	$t1, $t1, 1
memory[123] <= 32'h08000061;	//				j	sadouterloop
memory[124] <= 32'h11160002;	//	sadouterloopend:	beq	$t0, $s6, lteqcurrmin
memory[125] <= 32'h0116482a;	//				slt	$t1, $t0, $s6
memory[126] <= 32'h11200003;	//				beq	$t1, $0, lteqcurrminend
memory[127] <= 32'h0100b020;	//	lteqcurrmin:		add	$s6, $t0, $0
memory[128] <= 32'h01c01020;	//				add	$v0, $t6, $0
memory[129] <= 32'h01e01820;	//				add	$v1, $t7, $0
memory[130] <= 32'h03e00008;	//	lteqcurrminend:		jr	$ra
memory[131] <= 32'h21ef0001;	//	rightsubroutine:	addi	$t7, $t7, 1
memory[132] <= 32'h03e00008;	//				jr	$ra
memory[133] <= 32'h21ce0001;	//	downleftsubroutine:	addi	$t6, $t6, 1
memory[134] <= 32'h21efffff;	//				addi	$t7, $t7, -1
memory[135] <= 32'h03e00008;	//				jr	$ra
memory[136] <= 32'h21ceffff;	//	uprightsubroutine:	addi	$t6, $t6, -1
memory[137] <= 32'h21ef0001;	//				addi	$t7, $t7, 1
memory[138] <= 32'h03e00008;	//				jr	$ra
memory[139] <= 32'h21ce0001;	//	downsubroutine:		addi	$t6, $t6, 1
memory[140] <= 32'h03e00008;	//				jr	$ra
memory[141] <= 32'h21ceffff;	//	upsubroutine:		addi	$t6, $t6, -1
memory[142] <= 32'h21ef0001;	//				addi	$t7, $t7, 1
memory[143] <= 32'h03e00008;	//				jr	$ra































//regular dp with all test cases required.
/*
memory[0] <= 32'h23bdfffc;	//	main:			addi	$sp, $sp, -4
memory[1] <= 32'hafbf0000;	//				sw	$ra, 0($sp)
memory[2] <= 32'h34044df0;	//				ori	$a0, $zero, 19952
memory[3] <= 32'h34054e00;	//				ori	$a1, $zero, 19968
memory[4] <= 32'h34065200;	//				ori	$a2, $zero, 20992
memory[5] <= 32'h0c00000a;	//				jal	vbsme
memory[6] <= 32'h0c000008;	//				jal	print_result
memory[7] <= 32'h08000007;	//	exit:			j	exit
memory[8] <= 32'h00000000;	//	print_result:		nop
memory[9] <= 32'h03e00008;	//				jr	$ra
memory[10] <= 32'h8c900000;	//	vbsme:			lw	$s0, 0($a0)
memory[11] <= 32'h8c910004;	//				lw	$s1, 4($a0)
memory[12] <= 32'h8c920008;	//				lw	$s2, 8($a0)
memory[13] <= 32'h8c93000c;	//				lw	$s3, 12($a0)
memory[14] <= 32'h340e0000;	//				ori	$t6, $zero, 0
memory[15] <= 32'h340f0000;	//				ori	$t7, $zero, 0
memory[16] <= 32'h02124022;	//				sub	$t0, $s0, $s2
memory[17] <= 32'h71114002;	//				mul	$t0, $t0, $s1
memory[18] <= 32'h02334822;	//				sub	$t1, $s1, $s3
memory[19] <= 32'h0109a820;	//				add	$s5, $t0, $t1
memory[20] <= 32'hafa80004;	//				sw	$t0, 4($sp)
memory[21] <= 32'h34020000;	//				ori	$v0, $zero, 0
memory[22] <= 32'h34030000;	//				ori	$v1, $zero, 0
memory[23] <= 32'h3416270f;	//				ori	$s6, $zero, 9999
memory[24] <= 32'h23bdfffc;	//				addi	$sp, $sp, -4
memory[25] <= 32'hafbf0000;	//				sw	$ra, 0($sp)
memory[26] <= 32'h0271402a;	//				slt	$t0, $s3, $s1
memory[27] <= 32'h0250482a;	//				slt	$t1, $s2, $s0
memory[28] <= 32'h01094025;	//				or	$t0, $t0, $t1
memory[29] <= 32'h1100003c;	//				beq	$t0, $0, endzigzag
memory[30] <= 32'h0c00005e;	//				jal	sad
memory[31] <= 32'h02334022;	//				sub	$t0, $s1, $s3
memory[32] <= 32'h01e8402a;	//				slt	$t0, $t7, $t0
memory[33] <= 32'h11000002;	//				beq	$t0, $0, errordetectnexta
memory[34] <= 32'h0c000083;	//				jal	rightsubroutine
memory[35] <= 32'h08000028;	//				j	doneerrordetectright
memory[36] <= 32'h02124022;	//	errordetectnexta:	sub	$t0, $s0, $s2
memory[37] <= 32'h01c8402a;	//				slt	$t0, $t6, $t0
memory[38] <= 32'h11000033;	//				beq	$t0, $0, endzigzag
memory[39] <= 32'h0c00008b;	//				jal	downsubroutine
memory[40] <= 32'h0c00005e;	//	doneerrordetectright:	jal	sad
memory[41] <= 32'h71d14002;	//	zigzagloop:		mul	$t0, $t6, $s1
memory[42] <= 32'h010f4020;	//				add	$t0, $t0, $t7
memory[43] <= 32'h0115402a;	//				slt	$t0, $t0, $s5
memory[44] <= 32'h1100002d;	//				beq	$t0, $0, endzigzag
memory[45] <= 32'h20140001;	//				addi	$s4, $0, 1
memory[46] <= 32'h1280000e;	//	dlcollisiondetect:	beq	$s4, $0, edlcollisiondetect
memory[47] <= 32'h02124022;	//				sub	$t0, $s0, $s2
memory[48] <= 32'h01c8402a;	//				slt	$t0, $t6, $t0
memory[49] <= 32'h11000007;	//				beq	$t0, $0, downcollisiona
memory[50] <= 32'h000f402a;	//				slt	$t0, $0, $t7
memory[51] <= 32'h11000002;	//				beq	$t0, $0, leftcollisiona
memory[52] <= 32'h0c000085;	//				jal	downleftsubroutine
memory[53] <= 32'h0800003b;	//				j	downcollisionaend
memory[54] <= 32'h0c00008b;	//	leftcollisiona:		jal	downsubroutine
memory[55] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[56] <= 32'h0800003b;	//				j	downcollisionaend
memory[57] <= 32'h0c000083;	//	downcollisiona:		jal	rightsubroutine
memory[58] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[59] <= 32'h0c00005e;	//	downcollisionaend:	jal	sad
memory[60] <= 32'h0800002e;	//				j	dlcollisiondetect
memory[61] <= 32'h0c00005e;	//	edlcollisiondetect:	jal	sad
memory[62] <= 32'h71d14002;	//				mul	$t0, $t6, $s1
memory[63] <= 32'h010f4020;	//				add	$t0, $t0, $t7
memory[64] <= 32'h0115402a;	//				slt	$t0, $t0, $s5
memory[65] <= 32'h11000018;	//				beq	$t0, $0, endzigzag
memory[66] <= 32'h20140001;	//				addi	$s4, $0, 1
memory[67] <= 32'h12800014;	//	urcollisiondetect:	beq	$s4, $0, eurcollisiondetect
memory[68] <= 32'h000e402a;	//				slt	$t0, $0, $t6
memory[69] <= 32'h11000008;	//				beq	$t0, $0, upcollisiona
memory[70] <= 32'h02334022;	//				sub	$t0, $s1, $s3
memory[71] <= 32'h01e8402a;	//				slt	$t0, $t7, $t0
memory[72] <= 32'h11000002;	//				beq	$t0, $0, rightcollisiona
memory[73] <= 32'h0c000088;	//				jal	uprightsubroutine
memory[74] <= 32'h08000056;	//				j	upcollisionaend
memory[75] <= 32'h0c00008b;	//	rightcollisiona:	jal	downsubroutine
memory[76] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[77] <= 32'h08000056;	//				j	upcollisionaend
memory[78] <= 32'h02334022;	//	upcollisiona:		sub	$t0, $s1, $s3
memory[79] <= 32'h01e8402a;	//				slt	$t0, $t7, $t0
memory[80] <= 32'h11000003;	//				beq	$t0, $0, rightcollisionb
memory[81] <= 32'h0c000083;	//				jal	rightsubroutine
memory[82] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[83] <= 32'h08000056;	//				j	upcollisionaend
memory[84] <= 32'h0c00008b;	//	rightcollisionb:	jal	downsubroutine
memory[85] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[86] <= 32'h0c00005e;	//	upcollisionaend:	jal	sad
memory[87] <= 32'h08000043;	//				j	urcollisiondetect
memory[88] <= 32'h0c00005e;	//	eurcollisiondetect:	jal	sad
memory[89] <= 32'h08000029;	//				j	zigzagloop
memory[90] <= 32'h8fbf0000;	//	endzigzag:		lw	$ra, 0($sp)
memory[91] <= 32'h00000000;	//				nop
memory[92] <= 32'h00000000;	//				nop
memory[93] <= 32'h03e00008;	//				jr	$ra
memory[94] <= 32'h00000000;	//	sad:			nop
memory[95] <= 32'h00004020;	//				add	$t0, $0, $0
memory[96] <= 32'h00004820;	//				add	$t1, $0, $0
memory[97] <= 32'h0132582a;	//	sadouterloop:		slt	$t3, $t1, $s2
memory[98] <= 32'h11600019;	//				beq	$t3, $0, sadouterloopend
memory[99] <= 32'h00005020;	//				add	$t2, $0, $0
memory[100] <= 32'h0153582a;	//	sadinnerloop:		slt	$t3, $t2, $s3
memory[101] <= 32'h11600014;	//				beq	$t3, $0, sadinnerloopend
memory[102] <= 32'h012e5820;	//				add	$t3, $t1, $t6
memory[103] <= 32'h71715802;	//				mul	$t3, $t3, $s1
memory[104] <= 32'h016a5820;	//				add	$t3, $t3, $t2
memory[105] <= 32'h016f5820;	//				add	$t3, $t3, $t7
memory[106] <= 32'h000b5880;	//				sll	$t3, $t3, 2
memory[107] <= 32'h71336002;	//				mul	$t4, $t1, $s3
memory[108] <= 32'h018a6020;	//				add	$t4, $t4, $t2
memory[109] <= 32'h000c6080;	//				sll	$t4, $t4, 2
memory[110] <= 32'h00ab5820;	//				add	$t3, $a1, $t3
memory[111] <= 32'h00cc6020;	//				add	$t4, $a2, $t4
memory[112] <= 32'h8d6b0000;	//				lw	$t3, 0($t3)
memory[113] <= 32'h8d8c0000;	//				lw	$t4, 0($t4)
memory[114] <= 32'h016c5822;	//				sub	$t3, $t3, $t4
memory[115] <= 32'h0160602a;	//				slt	$t4, $t3, $0
memory[116] <= 32'h11800002;	//				beq	$t4, $0, absifend
memory[117] <= 32'h200dffff;	//				addi	$t5, $0, -1
memory[118] <= 32'h716d5802;	//				mul	$t3, $t3, $t5
memory[119] <= 32'h010b4020;	//	absifend:		add	$t0, $t0, $t3
memory[120] <= 32'h214a0001;	//				addi	$t2, $t2, 1
memory[121] <= 32'h08000064;	//				j	sadinnerloop
memory[122] <= 32'h21290001;	//	sadinnerloopend:	addi	$t1, $t1, 1
memory[123] <= 32'h08000061;	//				j	sadouterloop
memory[124] <= 32'h11160002;	//	sadouterloopend:	beq	$t0, $s6, lteqcurrmin
memory[125] <= 32'h0116482a;	//				slt	$t1, $t0, $s6
memory[126] <= 32'h11200003;	//				beq	$t1, $0, lteqcurrminend
memory[127] <= 32'h0100b020;	//	lteqcurrmin:		add	$s6, $t0, $0
memory[128] <= 32'h01c01020;	//				add	$v0, $t6, $0
memory[129] <= 32'h01e01820;	//				add	$v1, $t7, $0
memory[130] <= 32'h03e00008;	//	lteqcurrminend:		jr	$ra
memory[131] <= 32'h21ef0001;	//	rightsubroutine:	addi	$t7, $t7, 1
memory[132] <= 32'h03e00008;	//				jr	$ra
memory[133] <= 32'h21ce0001;	//	downleftsubroutine:	addi	$t6, $t6, 1
memory[134] <= 32'h21efffff;	//				addi	$t7, $t7, -1
memory[135] <= 32'h03e00008;	//				jr	$ra
memory[136] <= 32'h21ceffff;	//	uprightsubroutine:	addi	$t6, $t6, -1
memory[137] <= 32'h21ef0001;	//				addi	$t7, $t7, 1
memory[138] <= 32'h03e00008;	//				jr	$ra
memory[139] <= 32'h21ce0001;	//	downsubroutine:		addi	$t6, $t6, 1
memory[140] <= 32'h03e00008;	//				jr	$ra
memory[141] <= 32'h21ceffff;	//	upsubroutine:		addi	$t6, $t6, -1
memory[142] <= 32'h21ef0001;	//				addi	$t7, $t7, 1
memory[143] <= 32'h03e00008;	//				jr	$ra
*/


/*
 *  working vbsme code
 */

/*
memory[0] <= 32'h23bdfffc;	//	main:			addi	$sp, $sp, -4
memory[1] <= 32'hafbf0000;	//				sw	$ra, 0($sp)
memory[2] <= 32'h34044df0;	//				ori	$a0, $zero, 19952
memory[3] <= 32'h34054e00;	//				ori	$a1, $zero, 19968
memory[4] <= 32'h34065200;	//				ori	$a2, $zero, 20992
memory[5] <= 32'h0c00000a;	//				jal	vbsme
memory[6] <= 32'h0c000008;	//				jal	print_result
memory[7] <= 32'h08000007;	//	exit:			j	exit
memory[8] <= 32'h00000000;	//	print_result:		nop
memory[9] <= 32'h03e00008;	//				jr	$ra
memory[10] <= 32'h8c900000;	//	vbsme:			lw	$s0, 0($a0)
memory[11] <= 32'h8c910004;	//				lw	$s1, 4($a0)
memory[12] <= 32'h8c920008;	//				lw	$s2, 8($a0)
memory[13] <= 32'h8c93000c;	//				lw	$s3, 12($a0)
memory[14] <= 32'h340e0000;	//				ori	$t6, $zero, 0
memory[15] <= 32'h340f0000;	//				ori	$t7, $zero, 0
memory[16] <= 32'h02124022;	//				sub	$t0, $s0, $s2
memory[17] <= 32'h71114002;	//				mul	$t0, $t0, $s1
memory[18] <= 32'h02334822;	//				sub	$t1, $s1, $s3
memory[19] <= 32'h0109a820;	//				add	$s5, $t0, $t1
memory[20] <= 32'hafa80004;	//				sw	$t0, 4($sp)
memory[21] <= 32'h34020000;	//				ori	$v0, $zero, 0
memory[22] <= 32'h34030000;	//				ori	$v1, $zero, 0
memory[23] <= 32'h3416270f;	//				ori	$s6, $zero, 9999
memory[24] <= 32'h23bdfffc;	//				addi	$sp, $sp, -4
memory[25] <= 32'hafbf0000;	//				sw	$ra, 0($sp)
memory[26] <= 32'h0271402a;	//				slt	$t0, $s3, $s1
memory[27] <= 32'h0250482a;	//				slt	$t1, $s2, $s0
memory[28] <= 32'h01094025;	//				or	$t0, $t0, $t1
memory[29] <= 32'h11000047;	//				beq	$t0, $0, endzigzag
memory[30] <= 32'h0c00006b;	//				jal	sad
memory[31] <= 32'h02334022;	//				sub	$t0, $s1, $s3
memory[32] <= 32'h01e8402a;	//				slt	$t0, $t7, $t0
memory[33] <= 32'h11000002;	//				beq	$t0, $0, errordetectnexta
memory[34] <= 32'h0c0000f3;	//				jal	rightsubroutine
memory[35] <= 32'h08000028;	//				j	doneerrordetectright
memory[36] <= 32'h02124022;	//	errordetectnexta:	sub	$t0, $s0, $s2
memory[37] <= 32'h01c8402a;	//				slt	$t0, $t6, $t0
memory[38] <= 32'h1100003e;	//				beq	$t0, $0, endzigzag
memory[39] <= 32'h0c0000fd;	//				jal	downsubroutine
memory[40] <= 32'h0c00006b;	//	doneerrordetectright:	jal	sad
memory[41] <= 32'h00000000;	//	zigzagloop:		nop
memory[42] <= 32'h71d14002;	//				mul	$t0, $t6, $s1
memory[43] <= 32'h010f4020;	//				add	$t0, $t0, $t7
memory[44] <= 32'h0115402a;	//				slt	$t0, $t0, $s5
memory[45] <= 32'h11000037;	//				beq	$t0, $0, endzigzag
memory[46] <= 32'h20140001;	//				addi	$s4, $0, 1
memory[47] <= 32'h00000000;	//	dlcollisiondetect:	nop
memory[48] <= 32'h12800011;	//				beq	$s4, $0, edlcollisiondetect
memory[49] <= 32'h02124022;	//				sub	$t0, $s0, $s2
memory[50] <= 32'h01c8402a;	//				slt	$t0, $t6, $t0
memory[51] <= 32'h11000008;	//				beq	$t0, $0, downcollisiona
memory[52] <= 32'h000f402a;	//				slt	$t0, $0, $t7
memory[53] <= 32'h11000002;	//				beq	$t0, $0, leftcollisiona
memory[54] <= 32'h0c0000f6;	//				jal	downleftsubroutine
memory[55] <= 32'h0800003f;	//				j	downcollisionaend
memory[56] <= 32'h00000000;	//	leftcollisiona:		nop
memory[57] <= 32'h0c0000fd;	//				jal	downsubroutine
memory[58] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[59] <= 32'h0800003f;	//				j	downcollisionaend
memory[60] <= 32'h00000000;	//	downcollisiona:		nop
memory[61] <= 32'h0c0000f3;	//				jal	rightsubroutine
memory[62] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[63] <= 32'h00000000;	//	downcollisionaend:	nop
memory[64] <= 32'h0c00006b;	//				jal	sad
memory[65] <= 32'h0800002f;	//				j	dlcollisiondetect
memory[66] <= 32'h0c00006b;	//	edlcollisiondetect:	jal	sad
memory[67] <= 32'h71d14002;	//				mul	$t0, $t6, $s1
memory[68] <= 32'h010f4020;	//				add	$t0, $t0, $t7
memory[69] <= 32'h0115402a;	//				slt	$t0, $t0, $s5
memory[70] <= 32'h1100001e;	//				beq	$t0, $0, endzigzag
memory[71] <= 32'h20140001;	//				addi	$s4, $0, 1
memory[72] <= 32'h12800018;	//	urcollisiondetect:	beq	$s4, $0, eurcollisiondetect
memory[73] <= 32'h000e402a;	//				slt	$t0, $0, $t6
memory[74] <= 32'h11000009;	//				beq	$t0, $0, upcollisiona
memory[75] <= 32'h02334022;	//				sub	$t0, $s1, $s3
memory[76] <= 32'h01e8402a;	//				slt	$t0, $t7, $t0
memory[77] <= 32'h11000003;	//				beq	$t0, $0, rightcollisiona
memory[78] <= 32'h0c0000f9;	//				jal	uprightsubroutine
memory[79] <= 32'h00000000;	//				nop
memory[80] <= 32'h0800005d;	//				j	upcollisionaend
memory[81] <= 32'h0c0000fd;	//	rightcollisiona:	jal	downsubroutine
memory[82] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[83] <= 32'h0800005d;	//				j	upcollisionaend
memory[84] <= 32'h02334022;	//	upcollisiona:		sub	$t0, $s1, $s3
memory[85] <= 32'h01e8402a;	//				slt	$t0, $t7, $t0
memory[86] <= 32'h11000003;	//				beq	$t0, $0, rightcollisionb
memory[87] <= 32'h0c0000f3;	//				jal	rightsubroutine
memory[88] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[89] <= 32'h0800005d;	//				j	upcollisionaend
memory[90] <= 32'h00000000;	//	rightcollisionb:	nop
memory[91] <= 32'h0c0000fd;	//				jal	downsubroutine
memory[92] <= 32'h0000a020;	//				add	$s4, $0, $0
memory[93] <= 32'h00000000;	//	upcollisionaend:	nop
memory[94] <= 32'h0c00006b;	//				jal	sad
memory[95] <= 32'h00000000;	//				nop
memory[96] <= 32'h08000048;	//				j	urcollisiondetect
memory[97] <= 32'h00000000;	//	eurcollisiondetect:	nop
memory[98] <= 32'h0c00006b;	//				jal	sad
memory[99] <= 32'h00000000;	//				nop
memory[100] <= 32'h08000029;	//				j	zigzagloop
memory[101] <= 32'h00000000;	//	endzigzag:		nop
memory[102] <= 32'h00000000;	//				nop
memory[103] <= 32'h8fbf0000;	//				lw	$ra, 0($sp)
memory[104] <= 32'h00000000;	//				nop
memory[105] <= 32'h00000000;	//				nop
memory[106] <= 32'h03e00008;	//				jr	$ra
memory[107] <= 32'h00000000;	//	sad:			nop
memory[108] <= 32'h00000000;	//				nop
memory[109] <= 32'h00000000;	//				nop
memory[110] <= 32'h00000000;	//				nop
memory[111] <= 32'h00004020;	//				add	$t0, $0, $0
memory[112] <= 32'h00004820;	//				add	$t1, $0, $0
memory[113] <= 32'h00000000;	//	sadouterloop:		nop
memory[114] <= 32'h00000000;	//				nop
memory[115] <= 32'h00000000;	//				nop
memory[116] <= 32'h00000000;	//				nop
memory[117] <= 32'h0132582a;	//				slt	$t3, $t1, $s2
memory[118] <= 32'h00000000;	//				nop
memory[119] <= 32'h00000000;	//				nop
memory[120] <= 32'h00000000;	//				nop
memory[121] <= 32'h00000000;	//				nop
memory[122] <= 32'h11600065;	//				beq	$t3, $0, sadouterloopend
memory[123] <= 32'h00000000;	//				nop
memory[124] <= 32'h00000000;	//				nop
memory[125] <= 32'h00000000;	//				nop
memory[126] <= 32'h00000000;	//				nop
memory[127] <= 32'h00005020;	//				add	$t2, $0, $0
memory[128] <= 32'h00000000;	//	sadinnerloop:		nop
memory[129] <= 32'h00000000;	//				nop
memory[130] <= 32'h00000000;	//				nop
memory[131] <= 32'h00000000;	//				nop
memory[132] <= 32'h0153582a;	//				slt	$t3, $t2, $s3
memory[133] <= 32'h00000000;	//				nop
memory[134] <= 32'h00000000;	//				nop
memory[135] <= 32'h1160004e;	//				beq	$t3, $0, sadinnerloopend
memory[136] <= 32'h00000000;	//				nop
memory[137] <= 32'h00000000;	//				nop
memory[138] <= 32'h00000000;	//				nop
memory[139] <= 32'h00000000;	//				nop
memory[140] <= 32'h012e5820;	//				add	$t3, $t1, $t6
memory[141] <= 32'h00000000;	//				nop
memory[142] <= 32'h00000000;	//				nop
memory[143] <= 32'h00000000;	//				nop
memory[144] <= 32'h71715802;	//				mul	$t3, $t3, $s1
memory[145] <= 32'h00000000;	//				nop
memory[146] <= 32'h00000000;	//				nop
memory[147] <= 32'h00000000;	//				nop
memory[148] <= 32'h016a5820;	//				add	$t3, $t3, $t2
memory[149] <= 32'h00000000;	//				nop
memory[150] <= 32'h00000000;	//				nop
memory[151] <= 32'h00000000;	//				nop
memory[152] <= 32'h016f5820;	//				add	$t3, $t3, $t7
memory[153] <= 32'h00000000;	//				nop
memory[154] <= 32'h00000000;	//				nop
memory[155] <= 32'h00000000;	//				nop
memory[156] <= 32'h000b5880;	//				sll	$t3, $t3, 2
memory[157] <= 32'h00000000;	//				nop
memory[158] <= 32'h00000000;	//				nop
memory[159] <= 32'h00000000;	//				nop
memory[160] <= 32'h71336002;	//				mul	$t4, $t1, $s3
memory[161] <= 32'h00000000;	//				nop
memory[162] <= 32'h00000000;	//				nop
memory[163] <= 32'h00000000;	//				nop
memory[164] <= 32'h018a6020;	//				add	$t4, $t4, $t2
memory[165] <= 32'h00000000;	//				nop
memory[166] <= 32'h00000000;	//				nop
memory[167] <= 32'h00000000;	//				nop
memory[168] <= 32'h000c6080;	//				sll	$t4, $t4, 2
memory[169] <= 32'h00000000;	//				nop
memory[170] <= 32'h00000000;	//				nop
memory[171] <= 32'h00000000;	//				nop
memory[172] <= 32'h00ab5820;	//				add	$t3, $a1, $t3
memory[173] <= 32'h00000000;	//				nop
memory[174] <= 32'h00000000;	//				nop
memory[175] <= 32'h00000000;	//				nop
memory[176] <= 32'h00cc6020;	//				add	$t4, $a2, $t4
memory[177] <= 32'h00000000;	//				nop
memory[178] <= 32'h00000000;	//				nop
memory[179] <= 32'h00000000;	//				nop
memory[180] <= 32'h00000000;	//				nop
memory[181] <= 32'h8d6b0000;	//				lw	$t3, 0($t3)
memory[182] <= 32'h00000000;	//				nop
memory[183] <= 32'h00000000;	//				nop
memory[184] <= 32'h00000000;	//				nop
memory[185] <= 32'h00000000;	//				nop
memory[186] <= 32'h8d8c0000;	//				lw	$t4, 0($t4)
memory[187] <= 32'h00000000;	//				nop
memory[188] <= 32'h00000000;	//				nop
memory[189] <= 32'h00000000;	//				nop
memory[190] <= 32'h00000000;	//				nop
memory[191] <= 32'h016c5822;	//				sub	$t3, $t3, $t4
memory[192] <= 32'h00000000;	//				nop
memory[193] <= 32'h00000000;	//				nop
memory[194] <= 32'h00000000;	//				nop
memory[195] <= 32'h0160602a;	//				slt	$t4, $t3, $0
memory[196] <= 32'h00000000;	//				nop
memory[197] <= 32'h00000000;	//				nop
memory[198] <= 32'h00000000;	//				nop
memory[199] <= 32'h00000000;	//				nop
memory[200] <= 32'h11800002;	//				beq	$t4, $0, absifend
memory[201] <= 32'h200dffff;	//				addi	$t5, $0, -1
memory[202] <= 32'h716d5802;	//				mul	$t3, $t3, $t5
memory[203] <= 32'h00000000;	//	absifend:		nop
memory[204] <= 32'h00000000;	//				nop
memory[205] <= 32'h00000000;	//				nop
memory[206] <= 32'h00000000;	//				nop
memory[207] <= 32'h010b4020;	//				add	$t0, $t0, $t3
memory[208] <= 32'h214a0001;	//				addi	$t2, $t2, 1
memory[209] <= 32'h00000000;	//				nop
memory[210] <= 32'h00000000;	//				nop
memory[211] <= 32'h00000000;	//				nop
memory[212] <= 32'h00000000;	//				nop
memory[213] <= 32'h08000080;	//				j	sadinnerloop
memory[214] <= 32'h00000000;	//	sadinnerloopend:	nop
memory[215] <= 32'h00000000;	//				nop
memory[216] <= 32'h00000000;	//				nop
memory[217] <= 32'h00000000;	//				nop
memory[218] <= 32'h21290001;	//				addi	$t1, $t1, 1
memory[219] <= 32'h00000000;	//				nop
memory[220] <= 32'h00000000;	//				nop
memory[221] <= 32'h00000000;	//				nop
memory[222] <= 32'h00000000;	//				nop
memory[223] <= 32'h08000071;	//				j	sadouterloop
memory[224] <= 32'h00000000;	//	sadouterloopend:	nop
memory[225] <= 32'h00000000;	//				nop
memory[226] <= 32'h00000000;	//				nop
memory[227] <= 32'h00000000;	//				nop
memory[228] <= 32'h11160006;	//				beq	$t0, $s6, lteqcurrmin
memory[229] <= 32'h0116482a;	//				slt	$t1, $t0, $s6
memory[230] <= 32'h00000000;	//				nop
memory[231] <= 32'h00000000;	//				nop
memory[232] <= 32'h00000000;	//				nop
memory[233] <= 32'h00000000;	//				nop
memory[234] <= 32'h11200003;	//				beq	$t1, $0, lteqcurrminend
memory[235] <= 32'h0100b020;	//	lteqcurrmin:		add	$s6, $t0, $0
memory[236] <= 32'h01c01020;	//				add	$v0, $t6, $0
memory[237] <= 32'h01e01820;	//				add	$v1, $t7, $0
memory[238] <= 32'h00000000;	//	lteqcurrminend:		nop
memory[239] <= 32'h00000000;	//				nop
memory[240] <= 32'h00000000;	//				nop
memory[241] <= 32'h00000000;	//				nop
memory[242] <= 32'h03e00008;	//				jr	$ra
memory[243] <= 32'h00000000;	//	rightsubroutine:	nop
memory[244] <= 32'h21ef0001;	//				addi	$t7, $t7, 1
memory[245] <= 32'h03e00008;	//				jr	$ra
memory[246] <= 32'h21ce0001;	//	downleftsubroutine:	addi	$t6, $t6, 1
memory[247] <= 32'h21efffff;	//				addi	$t7, $t7, -1
memory[248] <= 32'h03e00008;	//				jr	$ra
memory[249] <= 32'h00000000;	//	uprightsubroutine:	nop
memory[250] <= 32'h21ceffff;	//				addi	$t6, $t6, -1
memory[251] <= 32'h21ef0001;	//				addi	$t7, $t7, 1
memory[252] <= 32'h03e00008;	//				jr	$ra
memory[253] <= 32'h21ce0001;	//	downsubroutine:		addi	$t6, $t6, 1
memory[254] <= 32'h03e00008;	//				jr	$ra
memory[255] <= 32'h21ceffff;	//	upsubroutine:		addi	$t6, $t6, -1
memory[256] <= 32'h21ef0001;	//				addi	$t7, $t7, 1
memory[257] <= 32'h03e00008;	//				jr	$ra
*/
















        //$readmemh("/home/mitch/Instruction_memory.txt", memory);
        
       /*
        //test case 9-14
        memory[0] <= 32'h20100001;	//	main:	addi	$s0, $zero, 1
        memory[1] <= 32'h20110001;    //        addi    $s1, $zero, 1
        memory[2] <= 32'h02118024;    //        and    $s0, $s0, $s1
        memory[3] <= 32'h02008024;    //        and    $s0, $s0, $zero
        memory[4] <= 32'h02308022;    //        sub    $s0, $s1, $s0
        memory[5] <= 32'h02008027;    //        nor    $s0, $s0, $zero
        memory[6] <= 32'h02008027;    //        nor    $s0, $s0, $zero
        memory[7] <= 32'h00008025;    //        or    $s0, $zero, $zero
        memory[8] <= 32'h02208025;    //        or    $s0, $s1, $zero
        memory[9] <= 32'h00108080;    //        sll    $s0, $s0, 2
        memory[10] <= 32'h02308004;    //        sllv    $s0, $s0, $s1
        memory[11] <= 32'h0200802a;    //        slt    $s0, $s0, $zero
        memory[12] <= 32'h0211802a;    //        slt    $s0, $s0, $s1
        memory[13] <= 32'h00118043;    //        sra    $s0, $s1, 1
        memory[14] <= 32'h00118007;    //        srav    $s0, $s1, $zero
        memory[15] <= 32'h00118042;    //        srl    $s0, $s1, 1
        memory[16] <= 32'h001180c0;    //        sll    $s0, $s1, 3
        memory[17] <= 32'h001080c2;    //        srl    $s0, $s0, 3
        memory[18] <= 32'h02308004;    //        sllv    $s0, $s0, $s1
        memory[19] <= 32'h02308006;    //        srlv    $s0, $s0, $s1
        memory[20] <= 32'h02118026;    //        xor    $s0, $s0, $s1
        memory[21] <= 32'h02118026;    //        xor    $s0, $s0, $s1
        memory[22] <= 32'h20120004;    //        addi    $s2, $zero, 4
        memory[23] <= 32'h72128002;    //        mul    $s0, $s0, $s2
        memory[24] <= 32'h22100004;    //        addi    $s0, $s0, 4
        memory[25] <= 32'h32100000;    //        andi    $s0, $s0, 0
        memory[26] <= 32'h36100001;    //        ori    $s0, $s0, 1
        memory[27] <= 32'h2a100000;    //        slti    $s0, $s0, 0
        memory[28] <= 32'h2a100001;    //        slti    $s0, $s0, 1
        memory[29] <= 32'h3a100001;    //        xori    $s0, $s0, 1
        memory[30] <= 32'h3a100001;    //        xori    $s0, $s0, 1
        memory[31] <= 32'h2010fffe;    //        addi    $s0, $zero, -2
        memory[32] <= 32'h20110002;    //        addi    $s1, $zero, 2
        memory[33] <= 32'h0230902b;    //        sltu    $s2, $s1, $s0
        memory[34] <= 32'h2e30fffe;    //        sltiu    $s0, $s1, -2
        memory[35] <= 32'h0220800a;    //        movz    $s0, $s1, $zero
        memory[36] <= 32'h0011800b;    //        movn    $s0, $zero, $s1
        memory[37] <= 32'h02328020;    //        add    $s0, $s1, $s2
        memory[38] <= 32'h2010fffe;    //        addi    $s0, $zero, -2
        memory[39] <= 32'h02308821;    //        addu    $s1, $s1, $s0
        memory[40] <= 32'h2411ffff;    //        addiu    $s1, $zero, -1
        memory[41] <= 32'h20120020;    //        addi    $s2, $zero, 32
        memory[42] <= 32'h02320018;    //        mult    $s1, $s2
        memory[43] <= 32'h0000a010;    //        mfhi    $s4
        memory[44] <= 32'h0000a812;    //        mflo    $s5
        memory[45] <= 32'h02320019;    //        multu    $s1, $s2
        memory[46] <= 32'h0000a010;    //        mfhi    $s4
        memory[47] <= 32'h0000a812;    //        mflo    $s5
        memory[48] <= 32'h72320000;    //        madd    $s1, $s2
        memory[49] <= 32'h0000a010;    //        mfhi    $s4
        memory[50] <= 32'h0000a812;    //        mflo    $s5
        memory[51] <= 32'h02400011;    //        mthi    $s2
        memory[52] <= 32'h02200013;    //        mtlo    $s1
        memory[53] <= 32'h0000a010;    //        mfhi    $s4
        memory[54] <= 32'h0000a812;    //        mflo    $s5
        memory[55] <= 32'h3231ffff;    //        andi    $s1, $s1, 65535
        memory[56] <= 32'h72920004;    //        msub    $s4, $s2
        memory[57] <= 32'h0000a010;    //        mfhi    $s4
        memory[58] <= 32'h0000a812;    //        mflo    $s5
        memory[59] <= 32'h20120001;    //        addi    $s2, $zero, 1
        memory[60] <= 32'h00328fc2;    //        rotr    $s1, $s2, 31
        memory[61] <= 32'h2014001f;    //        addi    $s4, $zero, 31
        memory[62] <= 32'h02918846;    //        rotrv    $s1, $s1, $s4
        memory[63] <= 32'h34110ff0;    //        ori    $s1, $zero, 0x0FF0
        memory[64] <= 32'h7c11a420;    //        seb    $s4, $s1
        memory[65] <= 32'h7c11a620;    //        seh    $s4, $s1
    */
        
        
        
        /*
memory[0] <= 32'h20100001;	//	main:		addi	$s0, $0, 1
    memory[1] <= 32'h20110001;    //            addi    $s1, $0, 1
    memory[2] <= 32'h12300022;    //            beq    $s1, $s0, checkone
    memory[3] <= 32'h00000000;    //    testtwo:    nop
    memory[4] <= 32'h00000000;    //            nop
    memory[5] <= 32'h00000000;    //            nop
    memory[6] <= 32'h00000000;    //            nop
    memory[7] <= 32'h20110002;    //            addi    $s1, $0, 2
    memory[8] <= 32'h20120002;    //            addi    $s2, $0, 2
    memory[9] <= 32'h1232001d;    //            beq    $s1, $s2, checktwo
    memory[10] <= 32'h00000000;    //    testthree:    nop
    memory[11] <= 32'h00000000;    //            nop
    memory[12] <= 32'h00000000;    //            nop
    memory[13] <= 32'h00000000;    //            nop
    memory[14] <= 32'h20100003;    //            addi    $s0, $0, 3
    memory[15] <= 32'h20110003;    //            addi    $s1, $0, 3
    memory[16] <= 32'h02119020;    //            add    $s2, $s0, $s1
    memory[17] <= 32'h02119820;    //            add    $s3, $s0, $s1
    memory[18] <= 32'h12720016;    //            beq    $s3, $s2, checkthree
    memory[19] <= 32'h00000000;    //    testfour:    nop
    memory[20] <= 32'h00000000;    //            nop
    memory[21] <= 32'h00000000;    //            nop
    memory[22] <= 32'h00000000;    //            nop
    memory[23] <= 32'h20100004;    //            addi    $s0, $0, 4
    memory[24] <= 32'h20110004;    //            addi    $s1, $0, 4
    memory[25] <= 32'h02119820;    //            add    $s3, $s0, $s1
    memory[26] <= 32'h02119020;    //            add    $s2, $s0, $s1
    memory[27] <= 32'h1272000f;    //            beq    $s3, $s2, checkfour
    memory[28] <= 32'h00000000;    //    testfive:    nop
    memory[29] <= 32'h00000000;    //            nop
    memory[30] <= 32'h00000000;    //            nop
    memory[31] <= 32'h00000000;    //            nop
    memory[32] <= 32'h20100005;    //            addi    $s0, $0, 5
    memory[33] <= 32'hac100000;    //            sw    $s0, 0($0)
    memory[34] <= 32'h8c110000;    //            lw    $s1, 0($0)
    memory[35] <= 32'h12200009;    //            beq    $s1, $0, checkfive
    memory[36] <= 32'h08000024;    //    end:        j    end
    memory[37] <= 32'h20160001;    //    checkone:    addi    $s6, $0, 1
    memory[38] <= 32'h08000003;    //            j    testtwo
    memory[39] <= 32'h20160002;    //    checktwo:    addi    $s6, $0, 2
    memory[40] <= 32'h0800000a;    //            j    testthree
    memory[41] <= 32'h20160003;    //    checkthree:    addi    $s6, $0, 3
    memory[42] <= 32'h08000013;    //            j    testfour
    memory[43] <= 32'h20160004;    //    checkfour:    addi    $s6, $0, 4
    memory[44] <= 32'h0800001c;    //            j    testfive
    memory[45] <= 32'h20160005;    //    checkfive:    addi    $s6, $0, 5
    memory[46] <= 32'h08000024;    //            j    end
        */
        
        
        
        
 /*
        
          //public test case Final Phase1
  memory[0] <= 32'h34120000;  //      main:           ori     $s2, $zero, 0
  memory[1] <= 32'h8e520000;    //            lw    $s2, 0($s2)

  memory[2] <= 32'h34130000;    //            ori    $s3, $zero, 0
  memory[3] <= 32'h8e730004;    //            lw    $s3, 4($s3)
  
  
  memory[4] <= 32'h02538820;    //            add    $s1, $s2, $s3
  memory[5] <= 32'h0233a022;    //            sub    $s4, $s1, $s3
  memory[6] <= 32'h02348822;    //            sub    $s1, $s1, $s4
  memory[7] <= 32'h7233a002;    //            mul    $s4, $s1, $s3
  
  
  memory[8] <= 32'h0233a022;    //            sub    $s4, $s1, $s3
  memory[9] <= 32'h02538820;    //            add    $s1, $s2, $s3
  memory[10] <= 32'h7234b002;    //            mul    $s6, $s1, $s4
  memory[11] <= 32'h02968822;    //            sub    $s1, $s4, $s6
  memory[12] <= 32'h02568820;    //            add    $s1, $s2, $s6
  memory[13] <= 32'h3631aaaa;    //            ori    $s1, $s1, 43690
  memory[14] <= 32'h00118a80;    //            sll    $s1, $s1, 10
  memory[15] <= 32'h22350000;    //            addi    $s5, $s1, 0
  memory[16] <= 32'h22b70000;    //            addi    $s7, $s5, 0
  memory[17] <= 32'h34120018;    //            ori    $s2, $zero, 24
  memory[18] <= 32'h8e510000;    //            lw    $s1, 0($s2)
  memory[19] <= 32'h0235a022;    //            sub    $s4, $s1, $s5
  memory[20] <= 32'h0237b024;    //            and    $s6, $s1, $s7
  memory[21] <= 32'h0236b825;    //            or    $s7, $s1, $s6
  memory[22] <= 32'h02339022;    //            sub    $s2, $s1, $s3
  memory[23] <= 32'h02554024;    //            and    $t0, $s2, $s5
  memory[24] <= 32'h02d24825;    //            or    $t1, $s6, $s2
  memory[25] <= 32'h02525020;    //            add    $t2, $s2, $s2
  memory[26] <= 32'h34110000;    //            ori    $s1, $zero, 0
  memory[27] <= 32'hae290004;    //            sw    $t1, 4($s1)
  memory[28] <= 32'h8e2a0004;    //            lw    $t2, 4($s1)
  memory[29] <= 32'h02339022;    //            sub    $s2, $s1, $s3
  memory[30] <= 32'h02555825;    //            or    $t3, $s2, $s5
  memory[31] <= 32'h02526020;    //            add    $t4, $s2, $s2
  memory[32] <= 32'h02525025;    //            or    $t2, $s2, $s2
  memory[33] <= 32'h02eaa020;    //            add    $s4, $s7, $t2
  memory[34] <= 32'h34090000;    //            ori    $t1, $zero, 0
  memory[35] <= 32'h8d280000;    //            lw    $t0, 0($t1)
  memory[36] <= 32'h8d2a0004;    //            lw    $t2, 4($t1)
  memory[37] <= 32'had2a0000;    //            sw    $t2, 0($t1)
  memory[38] <= 32'had280004;    //            sw    $t0, 4($t1)
  memory[39] <= 32'h8d280000;    //            lw    $t0, 0($t1)
  memory[40] <= 32'h8d2a0004;    //            lw    $t2, 4($t1)
  
  //branchy boi
  memory[41] <= 32'h34040018;    //            ori    $a0, $zero, 24
  memory[42] <= 32'h0800002d;    //            j    start
  //memory[42] <= 32'h08100038;    //            j    start
  memory[43] <= 32'h2004ffff;    //            addi    $a0, $zero, -1
  memory[44] <= 32'h2004ffff;    //            addi    $a0, $zero, -1
  memory[45] <= 32'h8c900004;    //    start:        lw    $s0, 4($a0)
  memory[46] <= 32'hac900000;    //            sw    $s0, 0($a0)
  memory[47] <= 32'h06010003;    //    branch1:    bgez    $s0, branch2
  //memory[47] <= 32'h060100d8;    //    branch1:    bgez    $s0, branch2
  memory[48] <= 32'h22100001;    //            addi    $s0, $s0, 1
  memory[49] <= 32'h0601fffd;    //            bgez    $s0, branch1
  memory[50] <= 32'h0800003d;    //            j    error
  memory[51] <= 32'h2010ffff;    //    branch2:    addi    $s0, $zero, -1
  memory[52] <= 32'h06000003;    //            bltz    $s0, branch3
  memory[53] <= 32'h20100001;    //            addi    $s0, $zero, 1
  memory[54] <= 32'h1e00fffc;    //            bgtz    $s0, branch2
  memory[55] <= 32'h0800003d;    //            j    error
  memory[56] <= 32'h06000003;    //    branch3:    bltz    $s0, done
  memory[57] <= 32'h2010ffff;    //            addi    $s0, $zero, -1
  memory[58] <= 32'h0600fffd;    //            bltz    $s0, branch3
  memory[59] <= 32'h0800003d;    //            j    error
  memory[60] <= 32'h0800003c;    //    done:        j    done
  memory[61] <= 32'h0800003d;    //    error:        j    error
        */
        
       /*             
       *public test case 15-18 without NOPS
       *
       */
       
      /*
      
      memory[0] <= 32'h34040000;    //    main:        ori    $a0, $zero, 0
      memory[1] <= 32'h08000004;    //            j    start
      memory[2] <= 32'h2004000a;    //            addi    $a0, $zero, 10
      memory[3] <= 32'h2004000a;    //            addi    $a0, $zero, 10
      memory[4] <= 32'h8c900004;    //    start:        lw    $s0, 4($a0)
      memory[5] <= 32'h8c900008;    //            lw    $s0, 8($a0)
      memory[6] <= 32'hac900000;    //            sw    $s0, 0($a0)
      memory[7] <= 32'hac90000c;    //            sw    $s0, 12($a0)
      memory[8] <= 32'h8c910000;    //            lw    $s1, 0($a0)
      memory[9] <= 32'h8c92000c;    //            lw    $s2, 12($a0)
      memory[10] <= 32'h12000003;    //            beq    $s0, $zero, branch1
      memory[11] <= 32'h02008820;    //            add    $s1, $s0, $zero
      memory[12] <= 32'h12110001;    //            beq    $s0, $s1, branch1
      memory[13] <= 32'h08000035;    //            j    error
      memory[14] <= 32'h2010ffff;    //    branch1:    addi    $s0, $zero, -1
      memory[15] <= 32'h0601fff4;    //            bgez    $s0, start
      memory[16] <= 32'h22100001;    //            addi    $s0, $s0, 1
      memory[17] <= 32'h06010001;    //            bgez    $s0, branch2
      memory[18] <= 32'h08000035;    //            j    error
      memory[19] <= 32'h2010ffff;    //    branch2:    addi    $s0, $zero, -1
      memory[20] <= 32'h1e000003;    //            bgtz    $s0, branch3
      memory[21] <= 32'h20100001;    //            addi    $s0, $zero, 1
      memory[22] <= 32'h1e000001;    //            bgtz    $s0, branch3
      memory[23] <= 32'h08000035;    //            j    error
      memory[24] <= 32'h06000003;    //    branch3:    bltz    $s0, branch4
      memory[25] <= 32'h2010ffff;    //            addi    $s0, $zero, -1
      memory[26] <= 32'h06000001;    //            bltz    $s0, branch4
      memory[27] <= 32'h08000035;    //            j    error
      memory[28] <= 32'h2011ffff;    //    branch4:    addi    $s1, $zero, -1
      memory[29] <= 32'h16110002;    //            bne    $s0, $s1, branch5
      memory[30] <= 32'h16000001;    //            bne    $s0, $zero, branch5
      memory[31] <= 32'h08000035;    //            j    error
      memory[32] <= 32'h20100080;    //    branch5:    addi    $s0, $zero, 128
      memory[33] <= 32'ha0900000;    //            sb    $s0, 0($a0)
      memory[34] <= 32'h80900000;    //            lb    $s0, 0($a0)
      memory[35] <= 32'h1a000001;    //            blez    $s0, branch6
      memory[36] <= 32'h08000035;    //            j    error
      memory[37] <= 32'h2010ffff;    //    branch6:    addi    $s0, $zero, -1
      memory[38] <= 32'ha4900000;    //            sh    $s0, 0($a0)
      memory[39] <= 32'h20100000;    //            addi    $s0, $zero, 0
      memory[40] <= 32'h84900000;    //            lh    $s0, 0($a0)
      memory[41] <= 32'h1a000001;    //            blez    $s0, branch7
      memory[42] <= 32'h08000035;    //            j    error
      memory[43] <= 32'h2010ffff;    //    branch7:    addi    $s0, $zero, -1
      memory[44] <= 32'h3c100001;    //            lui    $s0, 1
      memory[45] <= 32'h06010001;    //            bgez    $s0, branch8
      memory[46] <= 32'h08000035;    //            j    error
      memory[47] <= 32'h08000031;    //    branch8:    j    jump1
      memory[48] <= 32'h2210fffe;    //            addi    $s0, $s0, -2
      memory[49] <= 32'h0c000033;    //    jump1:        jal    jal1
      memory[50] <= 32'h08000004;    //            j    start
      memory[51] <= 32'h03e00008;    //    jal1:        jr    $ra
      memory[52] <= 32'h08000035;    //            j    error
      memory[53] <= 32'h00000008;    //    error:        jr    $zero
      memory[54] <= 32'h3402000a;    //            ori    $v0, $zero, 10
      memory[55] <= 32'h00000000;    //            nop
    */
  
        
        /*
        memory[0] <= 32'h08000009;    //   	 j    main
        memory[1] <= 32'h22100006;    //    tomato:    addi    $s0, $s0, 6
        memory[2] <= 32'h03e00008;    //   	 jr    $ra
        memory[3] <= 32'h22110005;    //    orange:    addi    $s1, $s0, 5
        memory[4] <= 32'h22120005;    //   	 addi    $s2, $s0, 5
        memory[5] <= 32'h22130005;    //   	 addi    $s3, $s0, 5
        memory[6] <= 32'h22140005;    //   	 addi    $s4, $s0, 5
        memory[7] <= 32'h22150005;    //   	 addi    $s5, $s0, 5
        memory[8] <= 32'h03e00008;    //   	 jr    $ra
        memory[9] <= 32'h34100004;    //    main:    ori    $s0, $zero, 4
        memory[10] <= 32'h0c000001;    //   	 jal    tomato
        memory[11] <= 32'h02108820;    //   	 add    $s1, $s0, $s0
        memory[12] <= 32'h02309020;    //   	 add    $s2, $s1, $s0
        memory[13] <= 32'h0c000003;    //   	 jal    orange
        */


        /*
         *
         *
         */
         
        /*
   memory[0] <= 32'h23bdfffc;	//	main:			addi	$sp, $sp, -4
        memory[1] <= 32'hafbf0000;    //                sw    $ra, 0($sp)
        memory[2] <= 32'h34040000;    //                ori    $a0, $zero, 0
        memory[3] <= 32'h34050010;    //                ori    $a1, $zero, 16
        memory[4] <= 32'h34060050;    //                ori    $a2, $zero, 80
        memory[5] <= 32'h0c000071;    //                jal    vbsme
        memory[6] <= 32'h0c00006f;    //                jal    print_result
        memory[7] <= 32'h34040060;    //                ori    $a0, $zero, 96
        memory[8] <= 32'h34050070;    //                ori    $a1, $zero, 112
        memory[9] <= 32'h34060470;    //                ori    $a2, $zero, 1136
        memory[10] <= 32'h0c000071;    //                jal    vbsme
        memory[11] <= 32'h0c00006f;    //                jal    print_result
        memory[12] <= 32'h340404b0;    //                ori    $a0, $zero, 1200
        memory[13] <= 32'h340504c0;    //                ori    $a1, $zero, 1216
        memory[14] <= 32'h340608c0;    //                ori    $a2, $zero, 2240
        memory[15] <= 32'h0c000071;    //                jal    vbsme
        memory[16] <= 32'h0c00006f;    //                jal    print_result
        memory[17] <= 32'h34040940;    //                ori    $a0, $zero, 2368
        memory[18] <= 32'h34050950;    //                ori    $a1, $zero, 2384
        memory[19] <= 32'h34060d50;    //                ori    $a2, $zero, 3408
        memory[20] <= 32'h0c000071;    //                jal    vbsme
        memory[21] <= 32'h0c00006f;    //                jal    print_result
        memory[22] <= 32'h34040dd0;    //                ori    $a0, $zero, 3536
        memory[23] <= 32'h34050de0;    //                ori    $a1, $zero, 3552
        memory[24] <= 32'h340611e0;    //                ori    $a2, $zero, 4576
        memory[25] <= 32'h0c000071;    //                jal    vbsme
        memory[26] <= 32'h0c00006f;    //                jal    print_result
        memory[27] <= 32'h34041220;    //                ori    $a0, $zero, 4640
        memory[28] <= 32'h34051230;    //                ori    $a1, $zero, 4656
        memory[29] <= 32'h34062230;    //                ori    $a2, $zero, 8752
        memory[30] <= 32'h0c000071;    //                jal    vbsme
        memory[31] <= 32'h0c00006f;    //                jal    print_result
        memory[32] <= 32'h34042430;    //                ori    $a0, $zero, 9264
        memory[33] <= 32'h34052440;    //                ori    $a1, $zero, 9280
        memory[34] <= 32'h34063440;    //                ori    $a2, $zero, 13376
        memory[35] <= 32'h0c000071;    //                jal    vbsme
        memory[36] <= 32'h0c00006f;    //                jal    print_result
        memory[37] <= 32'h34043480;    //                ori    $a0, $zero, 13440
        memory[38] <= 32'h34053490;    //                ori    $a1, $zero, 13456
        memory[39] <= 32'h34064490;    //                ori    $a2, $zero, 17552
        memory[40] <= 32'h0c000071;    //                jal    vbsme
        memory[41] <= 32'h0c00006f;    //                jal    print_result
        memory[42] <= 32'h34044510;    //                ori    $a0, $zero, 17680
        memory[43] <= 32'h34054520;    //                ori    $a1, $zero, 17696
        memory[44] <= 32'h34064920;    //                ori    $a2, $zero, 18720
        memory[45] <= 32'h0c000071;    //                jal    vbsme
        memory[46] <= 32'h0c00006f;    //                jal    print_result
        memory[47] <= 32'h340449a0;    //                ori    $a0, $zero, 18848
        memory[48] <= 32'h340549b0;    //                ori    $a1, $zero, 18864
        memory[49] <= 32'h34064db0;    //                ori    $a2, $zero, 19888
        memory[50] <= 32'h0c000071;    //                jal    vbsme
        memory[51] <= 32'h0c00006f;    //                jal    print_result
        memory[52] <= 32'h34044df0;    //                ori    $a0, $zero, 19952
        memory[53] <= 32'h34054e00;    //                ori    $a1, $zero, 19968
        memory[54] <= 32'h34065200;    //                ori    $a2, $zero, 20992
        memory[55] <= 32'h0c000071;    //                jal    vbsme
        memory[56] <= 32'h0c00006f;    //                jal    print_result
        memory[57] <= 32'h34045300;    //                ori    $a0, $zero, 21248
        memory[58] <= 32'h34055310;    //                ori    $a1, $zero, 21264
        memory[59] <= 32'h34066310;    //                ori    $a2, $zero, 25360
        memory[60] <= 32'h0c000071;    //                jal    vbsme
        memory[61] <= 32'h0c00006f;    //                jal    print_result
        memory[62] <= 32'h34046710;    //                ori    $a0, $zero, 26384
        memory[63] <= 32'h34056720;    //                ori    $a1, $zero, 26400
        memory[64] <= 32'h34066b20;    //                ori    $a2, $zero, 27424
        memory[65] <= 32'h0c000071;    //                jal    vbsme
        memory[66] <= 32'h0c00006f;    //                jal    print_result
        memory[67] <= 32'h34046b60;    //                ori    $a0, $zero, 27488
        memory[68] <= 32'h34056b70;    //                ori    $a1, $zero, 27504
        memory[69] <= 32'h34067b70;    //                ori    $a2, $zero, 31600
        memory[70] <= 32'h0c000071;    //                jal    vbsme
        memory[71] <= 32'h0c00006f;    //                jal    print_result
        memory[72] <= 32'h34047bb0;    //                ori    $a0, $zero, 31664
        memory[73] <= 32'h34057bc0;    //                ori    $a1, $zero, 31680
        memory[74] <= 32'h34067c00;    //                ori    $a2, $zero, 31744
        memory[75] <= 32'h0c000071;    //                jal    vbsme
        memory[76] <= 32'h0c00006f;    //                jal    print_result
        memory[77] <= 32'h34047c40;    //                ori    $a0, $zero, 31808
        memory[78] <= 32'h34057c50;    //                ori    $a1, $zero, 31824
        memory[79] <= 32'h34067c90;    //                ori    $a2, $zero, 31888
        memory[80] <= 32'h0c000071;    //                jal    vbsme
        memory[81] <= 32'h0c00006f;    //                jal    print_result
        memory[82] <= 32'h34047cd8;    //                ori    $a0, $zero, 31960
        memory[83] <= 32'h34057ce8;    //                ori    $a1, $zero, 31976
        memory[84] <= 32'h34067d58;    //                ori    $a2, $zero, 32088
        memory[85] <= 32'h0c000071;    //                jal    vbsme
        memory[86] <= 32'h0c00006f;    //                jal    print_result
        memory[87] <= 32'h34047da0;    //                ori    $a0, $zero, 32160
        memory[88] <= 32'h34057db0;    //                ori    $a1, $zero, 32176
        memory[89] <= 32'h34067e00;    //                ori    $a2, $zero, 32256
        memory[90] <= 32'h0c000071;    //                jal    vbsme
        memory[91] <= 32'h0c00006f;    //                jal    print_result
        memory[92] <= 32'h34047e20;    //                ori    $a0, $zero, 32288
        memory[93] <= 32'h34057e30;    //                ori    $a1, $zero, 32304
        memory[94] <= 32'h34067e80;    //                ori    $a2, $zero, 32384
        memory[95] <= 32'h0c000071;    //                jal    vbsme
        memory[96] <= 32'h0c00006f;    //                jal    print_result
        memory[97] <= 32'h34047e8c;    //                ori    $a0, $zero, 32396
        memory[98] <= 32'h34057e9c;    //                ori    $a1, $zero, 32412
        memory[99] <= 32'h34067eec;    //                ori    $a2, $zero, 32492
        memory[100] <= 32'h0c000071;    //                jal    vbsme
        memory[101] <= 32'h0c00006f;    //                jal    print_result
        memory[102] <= 32'h34047ef8;    //                ori    $a0, $zero, 32504
        memory[103] <= 32'h34057f08;    //                ori    $a1, $zero, 32520
        memory[104] <= 32'h34067f50;    //                ori    $a2, $zero, 32592
        memory[105] <= 32'h0c000071;    //                jal    vbsme
        memory[106] <= 32'h0c00006f;    //                jal    print_result
        memory[107] <= 32'h8fbf0000;    //                lw    $ra, 0($sp)
        memory[108] <= 32'h23bd0004;    //                addi    $sp, $sp, 4
        memory[109] <= 32'h3402000a;    //    exit:            ori    $v0, $zero, 10
        memory[110] <= 32'h00000000;    //                nop
        memory[111] <= 32'h00000000;    //    print_result:        nop
        memory[112] <= 32'h03e00008;    //                jr    $ra
        memory[113] <= 32'h8c900000;    //    vbsme:            lw    $s0, 0($a0)
        memory[114] <= 32'h8c910004;    //                lw    $s1, 4($a0)
        memory[115] <= 32'h8c920008;    //                lw    $s2, 8($a0)
        memory[116] <= 32'h8c93000c;    //                lw    $s3, 12($a0)
        memory[117] <= 32'h340e0000;    //                ori    $t6, $zero, 0
        memory[118] <= 32'h340f0000;    //                ori    $t7, $zero, 0
        memory[119] <= 32'h02124022;    //                sub    $t0, $s0, $s2
        memory[120] <= 32'h71114002;    //                mul    $t0, $t0, $s1
        memory[121] <= 32'h02334822;    //                sub    $t1, $s1, $s3
        memory[122] <= 32'h0109a820;    //                add    $s5, $t0, $t1
        memory[123] <= 32'hafa80004;    //                sw    $t0, 4($sp)
        memory[124] <= 32'h34020000;    //                ori    $v0, $zero, 0
        memory[125] <= 32'h34030000;    //                ori    $v1, $zero, 0
        memory[126] <= 32'h3416270f;    //                ori    $s6, $zero, 9999
        memory[127] <= 32'h23bdfffc;    //                addi    $sp, $sp, -4
        memory[128] <= 32'hafbf0000;    //                sw    $ra, 0($sp)
        memory[129] <= 32'h0271402a;    //                slt    $t0, $s3, $s1
        memory[130] <= 32'h0250482a;    //                slt    $t1, $s2, $s0
        memory[131] <= 32'h01094025;    //                or    $t0, $t0, $t1
        memory[132] <= 32'h11000047;    //                beq    $t0, $0, endzigzag
        memory[133] <= 32'h0c0000d2;    //                jal    sad
        memory[134] <= 32'h02334022;    //                sub    $t0, $s1, $s3
        memory[135] <= 32'h01e8402a;    //                slt    $t0, $t7, $t0
        memory[136] <= 32'h11000002;    //                beq    $t0, $0, errordetectnexta
        memory[137] <= 32'h0c0000f8;    //                jal    rightsubroutine
        memory[138] <= 32'h0800008f;    //                j    doneerrordetectright
        memory[139] <= 32'h02124022;    //    errordetectnexta:    sub    $t0, $s0, $s2
        memory[140] <= 32'h01c8402a;    //                slt    $t0, $t6, $t0
        memory[141] <= 32'h1100003e;    //                beq    $t0, $0, endzigzag
        memory[142] <= 32'h0c000102;    //                jal    downsubroutine
        memory[143] <= 32'h0c0000d2;    //    doneerrordetectright:    jal    sad
        memory[144] <= 32'h00000000;    //    zigzagloop:        nop
        memory[145] <= 32'h71d14002;    //                mul    $t0, $t6, $s1
        memory[146] <= 32'h010f4020;    //                add    $t0, $t0, $t7
        memory[147] <= 32'h0115402a;    //                slt    $t0, $t0, $s5
        memory[148] <= 32'h11000037;    //                beq    $t0, $0, endzigzag
        memory[149] <= 32'h20140001;    //                addi    $s4, $0, 1
        memory[150] <= 32'h00000000;    //    dlcollisiondetect:    nop
        memory[151] <= 32'h12800011;    //                beq    $s4, $0, edlcollisiondetect
        memory[152] <= 32'h02124022;    //                sub    $t0, $s0, $s2
        memory[153] <= 32'h01c8402a;    //                slt    $t0, $t6, $t0
        memory[154] <= 32'h11000008;    //                beq    $t0, $0, downcollisiona
        memory[155] <= 32'h000f402a;    //                slt    $t0, $0, $t7
        memory[156] <= 32'h11000002;    //                beq    $t0, $0, leftcollisiona
        memory[157] <= 32'h0c0000fb;    //                jal    downleftsubroutine
        memory[158] <= 32'h080000a6;    //                j    downcollisionaend
        memory[159] <= 32'h00000000;    //    leftcollisiona:        nop
        memory[160] <= 32'h0c000102;    //                jal    downsubroutine
        memory[161] <= 32'h0000a020;    //                add    $s4, $0, $0
        memory[162] <= 32'h080000a6;    //                j    downcollisionaend
        memory[163] <= 32'h00000000;    //    downcollisiona:        nop
        memory[164] <= 32'h0c0000f8;    //                jal    rightsubroutine
        memory[165] <= 32'h0000a020;    //                add    $s4, $0, $0
        memory[166] <= 32'h00000000;    //    downcollisionaend:    nop
        memory[167] <= 32'h0c0000d2;    //                jal    sad
        memory[168] <= 32'h08000096;    //                j    dlcollisiondetect
        memory[169] <= 32'h0c0000d2;    //    edlcollisiondetect:    jal    sad
        memory[170] <= 32'h71d14002;    //                mul    $t0, $t6, $s1
        memory[171] <= 32'h010f4020;    //                add    $t0, $t0, $t7
        memory[172] <= 32'h0115402a;    //                slt    $t0, $t0, $s5
        memory[173] <= 32'h1100001e;    //                beq    $t0, $0, endzigzag
        memory[174] <= 32'h20140001;    //                addi    $s4, $0, 1
        memory[175] <= 32'h12800018;    //    urcollisiondetect:    beq    $s4, $0, eurcollisiondetect
        memory[176] <= 32'h000e402a;    //                slt    $t0, $0, $t6
        memory[177] <= 32'h11000009;    //                beq    $t0, $0, upcollisiona
        memory[178] <= 32'h02334022;    //                sub    $t0, $s1, $s3
        memory[179] <= 32'h01e8402a;    //                slt    $t0, $t7, $t0
        memory[180] <= 32'h11000003;    //                beq    $t0, $0, rightcollisiona
        memory[181] <= 32'h0c0000fe;    //                jal    uprightsubroutine
        memory[182] <= 32'h00000000;    //                nop
        memory[183] <= 32'h080000c4;    //                j    upcollisionaend
        memory[184] <= 32'h0c000102;    //    rightcollisiona:    jal    downsubroutine
        memory[185] <= 32'h0000a020;    //                add    $s4, $0, $0
        memory[186] <= 32'h080000c4;    //                j    upcollisionaend
        memory[187] <= 32'h02334022;    //    upcollisiona:        sub    $t0, $s1, $s3
        memory[188] <= 32'h01e8402a;    //                slt    $t0, $t7, $t0
        memory[189] <= 32'h11000003;    //                beq    $t0, $0, rightcollisionb
        memory[190] <= 32'h0c0000f8;    //                jal    rightsubroutine
        memory[191] <= 32'h0000a020;    //                add    $s4, $0, $0
        memory[192] <= 32'h080000c4;    //                j    upcollisionaend
        memory[193] <= 32'h00000000;    //    rightcollisionb:    nop
        memory[194] <= 32'h0c000102;    //                jal    downsubroutine
        memory[195] <= 32'h0000a020;    //                add    $s4, $0, $0
        memory[196] <= 32'h00000000;    //    upcollisionaend:    nop
        memory[197] <= 32'h0c0000d2;    //                jal    sad
        memory[198] <= 32'h00000000;    //                nop
        memory[199] <= 32'h080000af;    //                j    urcollisiondetect
        memory[200] <= 32'h00000000;    //    eurcollisiondetect:    nop
        memory[201] <= 32'h0c0000d2;    //                jal    sad
        memory[202] <= 32'h00000000;    //                nop
        memory[203] <= 32'h08000090;    //                j    zigzagloop
        memory[204] <= 32'h00000000;    //    endzigzag:        nop
        memory[205] <= 32'h00000000;    //                nop
        memory[206] <= 32'h8fbf0000;    //                lw    $ra, 0($sp)
        memory[207] <= 32'h00000000;    //                nop
        memory[208] <= 32'h00000000;    //                nop
        memory[209] <= 32'h03e00008;    //                jr    $ra
        memory[210] <= 32'h00004020;    //    sad:            add    $t0, $0, $0
        memory[211] <= 32'h00004820;    //                add    $t1, $0, $0
        memory[212] <= 32'h0132582a;    //    sadouterloop:        slt    $t3, $t1, $s2
        memory[213] <= 32'h1160001a;    //                beq    $t3, $0, sadouterloopend
        memory[214] <= 32'h00005020;    //                add    $t2, $0, $0
        memory[215] <= 32'h0153582a;    //    sadinnerloop:        slt    $t3, $t2, $s3
        memory[216] <= 32'h11600014;    //                beq    $t3, $0, sadinnerloopend
        memory[217] <= 32'h012e5820;    //                add    $t3, $t1, $t6
        memory[218] <= 32'h71715802;    //                mul    $t3, $t3, $s1
        memory[219] <= 32'h016a5820;    //                add    $t3, $t3, $t2
        memory[220] <= 32'h016f5820;    //                add    $t3, $t3, $t7
        memory[221] <= 32'h000b5880;    //                sll    $t3, $t3, 2
        memory[222] <= 32'h71336002;    //                mul    $t4, $t1, $s3
        memory[223] <= 32'h018a6020;    //                add    $t4, $t4, $t2
        memory[224] <= 32'h000c6080;    //                sll    $t4, $t4, 2
        memory[225] <= 32'h00ab5820;    //                add    $t3, $a1, $t3
        memory[226] <= 32'h00cc6020;    //                add    $t4, $a2, $t4
        memory[227] <= 32'h8d6b0000;    //                lw    $t3, 0($t3)
        memory[228] <= 32'h8d8c0000;    //                lw    $t4, 0($t4)
        memory[229] <= 32'h016c5822;    //                sub    $t3, $t3, $t4
        memory[230] <= 32'h0160602a;    //                slt    $t4, $t3, $0
        memory[231] <= 32'h11800002;    //                beq    $t4, $0, absifend
        memory[232] <= 32'h200dffff;    //                addi    $t5, $0, -1
        memory[233] <= 32'h716d5802;    //                mul    $t3, $t3, $t5
        memory[234] <= 32'h010b4020;    //    absifend:        add    $t0, $t0, $t3
        memory[235] <= 32'h214a0001;    //                addi    $t2, $t2, 1
        memory[236] <= 32'h080000d7;    //                j    sadinnerloop
        memory[237] <= 32'h00000000;    //    sadinnerloopend:    nop
        memory[238] <= 32'h21290001;    //                addi    $t1, $t1, 1
        memory[239] <= 32'h080000d4;    //                j    sadouterloop
        memory[240] <= 32'h11160002;    //    sadouterloopend:    beq    $t0, $s6, lteqcurrmin
        memory[241] <= 32'h0116482a;    //                slt    $t1, $t0, $s6
        memory[242] <= 32'h11200003;    //                beq    $t1, $0, lteqcurrminend
        memory[243] <= 32'h0100b020;    //    lteqcurrmin:        add    $s6, $t0, $0
        memory[244] <= 32'h01c01020;    //                add    $v0, $t6, $0
        memory[245] <= 32'h01e01820;    //                add    $v1, $t7, $0
        memory[246] <= 32'h00000000;    //    lteqcurrminend:        nop
        memory[247] <= 32'h03e00008;    //                jr    $ra
        memory[248] <= 32'h00000000;    //    rightsubroutine:    nop
        memory[249] <= 32'h21ef0001;    //                addi    $t7, $t7, 1
        memory[250] <= 32'h03e00008;    //                jr    $ra
        memory[251] <= 32'h21ce0001;    //    downleftsubroutine:    addi    $t6, $t6, 1
        memory[252] <= 32'h21efffff;    //                addi    $t7, $t7, -1
        memory[253] <= 32'h03e00008;    //                jr    $ra
        memory[254] <= 32'h00000000;    //    uprightsubroutine:    nop
        memory[255] <= 32'h21ceffff;    //                addi    $t6, $t6, -1
        memory[256] <= 32'h21ef0001;    //                addi    $t7, $t7, 1
        memory[257] <= 32'h03e00008;    //                jr    $ra
        memory[258] <= 32'h21ce0001;    //    downsubroutine:        addi    $t6, $t6, 1
        memory[259] <= 32'h03e00008;    //                jr    $ra
        memory[260] <= 32'h21ceffff;    //    upsubroutine:        addi    $t6, $t6, -1
        memory[261] <= 32'h21ef0001;    //                addi    $t7, $t7, 1
        memory[262] <= 32'h03e00008;    //                jr    $ra

*/



/*
    
    memory[0] <= 32'h23bdfffc;	//	main:			addi	$sp, $sp, -4
    memory[1] <= 32'h00000000;    //                nop
    memory[2] <= 32'h00000000;    //                nop
    memory[3] <= 32'h00000000;    //                nop
    memory[4] <= 32'h00000000;    //                nop
    memory[5] <= 32'hafbf0000;    //                sw    $ra, 0($sp)
    memory[6] <= 32'h00000000;    //                nop
    memory[7] <= 32'h00000000;    //                nop
    memory[8] <= 32'h00000000;    //                nop
    memory[9] <= 32'h00000000;    //                nop
    memory[10] <= 32'h34040000;    //                ori    $a0, $zero, 0
    memory[11] <= 32'h34050010;    //                ori    $a1, $zero, 16
    memory[12] <= 32'h34060050;    //                ori    $a2, $zero, 80
    memory[13] <= 32'h0c00017f;    //                jal    vbsme
    memory[14] <= 32'h00000000;    //                nop
    memory[15] <= 32'h00000000;    //                nop
    memory[16] <= 32'h00000000;    //                nop
    memory[17] <= 32'h00000000;    //                nop
    memory[18] <= 32'h0c00012f;    //                jal    print_result
    memory[19] <= 32'h00000000;    //                nop
    memory[20] <= 32'h00000000;    //                nop
    memory[21] <= 32'h00000000;    //                nop
    memory[22] <= 32'h00000000;    //                nop
    memory[23] <= 32'h34040060;    //                ori    $a0, $zero, 96
    memory[24] <= 32'h34050070;    //                ori    $a1, $zero, 112
    memory[25] <= 32'h34060470;    //                ori    $a2, $zero, 1136
    memory[26] <= 32'h0c00017f;    //                jal    vbsme
    memory[27] <= 32'h00000000;    //                nop
    memory[28] <= 32'h00000000;    //                nop
    memory[29] <= 32'h00000000;    //                nop
    memory[30] <= 32'h00000000;    //                nop
    memory[31] <= 32'h0c00012f;    //                jal    print_result
    memory[32] <= 32'h00000000;    //                nop
    memory[33] <= 32'h00000000;    //                nop
    memory[34] <= 32'h00000000;    //                nop
    memory[35] <= 32'h00000000;    //                nop
    memory[36] <= 32'h340404b0;    //                ori    $a0, $zero, 1200
    memory[37] <= 32'h340504c0;    //                ori    $a1, $zero, 1216
    memory[38] <= 32'h340608c0;    //                ori    $a2, $zero, 2240
    memory[39] <= 32'h0c00017f;    //                jal    vbsme
    memory[40] <= 32'h00000000;    //                nop
    memory[41] <= 32'h00000000;    //                nop
    memory[42] <= 32'h00000000;    //                nop
    memory[43] <= 32'h00000000;    //                nop
    memory[44] <= 32'h0c00012f;    //                jal    print_result
    memory[45] <= 32'h00000000;    //                nop
    memory[46] <= 32'h00000000;    //                nop
    memory[47] <= 32'h00000000;    //                nop
    memory[48] <= 32'h00000000;    //                nop
    memory[49] <= 32'h34040940;    //                ori    $a0, $zero, 2368
    memory[50] <= 32'h34050950;    //                ori    $a1, $zero, 2384
    memory[51] <= 32'h34060d50;    //                ori    $a2, $zero, 3408
    memory[52] <= 32'h0c00017f;    //                jal    vbsme
    memory[53] <= 32'h00000000;    //                nop
    memory[54] <= 32'h00000000;    //                nop
    memory[55] <= 32'h00000000;    //                nop
    memory[56] <= 32'h00000000;    //                nop
    memory[57] <= 32'h0c00012f;    //                jal    print_result
    memory[58] <= 32'h00000000;    //                nop
    memory[59] <= 32'h00000000;    //                nop
    memory[60] <= 32'h00000000;    //                nop
    memory[61] <= 32'h00000000;    //                nop
    memory[62] <= 32'h34040dd0;    //                ori    $a0, $zero, 3536
    memory[63] <= 32'h34050de0;    //                ori    $a1, $zero, 3552
    memory[64] <= 32'h340611e0;    //                ori    $a2, $zero, 4576
    memory[65] <= 32'h0c00017f;    //                jal    vbsme
    memory[66] <= 32'h00000000;    //                nop
    memory[67] <= 32'h00000000;    //                nop
    memory[68] <= 32'h00000000;    //                nop
    memory[69] <= 32'h00000000;    //                nop
    memory[70] <= 32'h0c00012f;    //                jal    print_result
    memory[71] <= 32'h00000000;    //                nop
    memory[72] <= 32'h00000000;    //                nop
    memory[73] <= 32'h00000000;    //                nop
    memory[74] <= 32'h00000000;    //                nop
    memory[75] <= 32'h34041220;    //                ori    $a0, $zero, 4640
    memory[76] <= 32'h34051230;    //                ori    $a1, $zero, 4656
    memory[77] <= 32'h34062230;    //                ori    $a2, $zero, 8752
    memory[78] <= 32'h0c00017f;    //                jal    vbsme
    memory[79] <= 32'h00000000;    //                nop
    memory[80] <= 32'h00000000;    //                nop
    memory[81] <= 32'h00000000;    //                nop
    memory[82] <= 32'h00000000;    //                nop
    memory[83] <= 32'h0c00012f;    //                jal    print_result
    memory[84] <= 32'h00000000;    //                nop
    memory[85] <= 32'h00000000;    //                nop
    memory[86] <= 32'h00000000;    //                nop
    memory[87] <= 32'h00000000;    //                nop
    memory[88] <= 32'h34042430;    //                ori    $a0, $zero, 9264
    memory[89] <= 32'h34052440;    //                ori    $a1, $zero, 9280
    memory[90] <= 32'h34063440;    //                ori    $a2, $zero, 13376
    memory[91] <= 32'h0c00017f;    //                jal    vbsme
    memory[92] <= 32'h00000000;    //                nop
    memory[93] <= 32'h00000000;    //                nop
    memory[94] <= 32'h00000000;    //                nop
    memory[95] <= 32'h00000000;    //                nop
    memory[96] <= 32'h0c00012f;    //                jal    print_result
    memory[97] <= 32'h00000000;    //                nop
    memory[98] <= 32'h00000000;    //                nop
    memory[99] <= 32'h00000000;    //                nop
    memory[100] <= 32'h00000000;    //                nop
    memory[101] <= 32'h34043480;    //                ori    $a0, $zero, 13440
    memory[102] <= 32'h34053490;    //                ori    $a1, $zero, 13456
    memory[103] <= 32'h34064490;    //                ori    $a2, $zero, 17552
    memory[104] <= 32'h0c00017f;    //                jal    vbsme
    memory[105] <= 32'h00000000;    //                nop
    memory[106] <= 32'h00000000;    //                nop
    memory[107] <= 32'h00000000;    //                nop
    memory[108] <= 32'h00000000;    //                nop
    memory[109] <= 32'h0c00012f;    //                jal    print_result
    memory[110] <= 32'h00000000;    //                nop
    memory[111] <= 32'h00000000;    //                nop
    memory[112] <= 32'h00000000;    //                nop
    memory[113] <= 32'h00000000;    //                nop
    memory[114] <= 32'h34044510;    //                ori    $a0, $zero, 17680
    memory[115] <= 32'h34054520;    //                ori    $a1, $zero, 17696
    memory[116] <= 32'h34064920;    //                ori    $a2, $zero, 18720
    memory[117] <= 32'h0c00017f;    //                jal    vbsme
    memory[118] <= 32'h00000000;    //                nop
    memory[119] <= 32'h00000000;    //                nop
    memory[120] <= 32'h00000000;    //                nop
    memory[121] <= 32'h00000000;    //                nop
    memory[122] <= 32'h0c00012f;    //                jal    print_result
    memory[123] <= 32'h00000000;    //                nop
    memory[124] <= 32'h00000000;    //                nop
    memory[125] <= 32'h00000000;    //                nop
    memory[126] <= 32'h00000000;    //                nop
    memory[127] <= 32'h340449a0;    //                ori    $a0, $zero, 18848
    memory[128] <= 32'h340549b0;    //                ori    $a1, $zero, 18864
    memory[129] <= 32'h34064db0;    //                ori    $a2, $zero, 19888
    memory[130] <= 32'h0c00017f;    //                jal    vbsme
    memory[131] <= 32'h00000000;    //                nop
    memory[132] <= 32'h00000000;    //                nop
    memory[133] <= 32'h00000000;    //                nop
    memory[134] <= 32'h00000000;    //                nop
    memory[135] <= 32'h0c00012f;    //                jal    print_result
    memory[136] <= 32'h00000000;    //                nop
    memory[137] <= 32'h00000000;    //                nop
    memory[138] <= 32'h00000000;    //                nop
    memory[139] <= 32'h00000000;    //                nop
    memory[140] <= 32'h34044df0;    //                ori    $a0, $zero, 19952
    memory[141] <= 32'h34054e00;    //                ori    $a1, $zero, 19968
    memory[142] <= 32'h34065200;    //                ori    $a2, $zero, 20992
    memory[143] <= 32'h0c00017f;    //                jal    vbsme
    memory[144] <= 32'h00000000;    //                nop
    memory[145] <= 32'h00000000;    //                nop
    memory[146] <= 32'h00000000;    //                nop
    memory[147] <= 32'h00000000;    //                nop
    memory[148] <= 32'h0c00012f;    //                jal    print_result
    memory[149] <= 32'h00000000;    //                nop
    memory[150] <= 32'h00000000;    //                nop
    memory[151] <= 32'h00000000;    //                nop
    memory[152] <= 32'h00000000;    //                nop
    memory[153] <= 32'h34045300;    //                ori    $a0, $zero, 21248
    memory[154] <= 32'h34055310;    //                ori    $a1, $zero, 21264
    memory[155] <= 32'h34066310;    //                ori    $a2, $zero, 25360
    memory[156] <= 32'h0c00017f;    //                jal    vbsme
    memory[157] <= 32'h00000000;    //                nop
    memory[158] <= 32'h00000000;    //                nop
    memory[159] <= 32'h00000000;    //                nop
    memory[160] <= 32'h00000000;    //                nop
    memory[161] <= 32'h0c00012f;    //                jal    print_result
    memory[162] <= 32'h00000000;    //                nop
    memory[163] <= 32'h00000000;    //                nop
    memory[164] <= 32'h00000000;    //                nop
    memory[165] <= 32'h00000000;    //                nop
    memory[166] <= 32'h34046710;    //                ori    $a0, $zero, 26384
    memory[167] <= 32'h34056720;    //                ori    $a1, $zero, 26400
    memory[168] <= 32'h34066b20;    //                ori    $a2, $zero, 27424
    memory[169] <= 32'h0c00017f;    //                jal    vbsme
    memory[170] <= 32'h00000000;    //                nop
    memory[171] <= 32'h00000000;    //                nop
    memory[172] <= 32'h00000000;    //                nop
    memory[173] <= 32'h00000000;    //                nop
    memory[174] <= 32'h0c00012f;    //                jal    print_result
    memory[175] <= 32'h00000000;    //                nop
    memory[176] <= 32'h00000000;    //                nop
    memory[177] <= 32'h00000000;    //                nop
    memory[178] <= 32'h00000000;    //                nop
    memory[179] <= 32'h34046b60;    //                ori    $a0, $zero, 27488
    memory[180] <= 32'h34056b70;    //                ori    $a1, $zero, 27504
    memory[181] <= 32'h34067b70;    //                ori    $a2, $zero, 31600
    memory[182] <= 32'h0c00017f;    //                jal    vbsme
    memory[183] <= 32'h00000000;    //                nop
    memory[184] <= 32'h00000000;    //                nop
    memory[185] <= 32'h00000000;    //                nop
    memory[186] <= 32'h00000000;    //                nop
    memory[187] <= 32'h0c00012f;    //                jal    print_result
    memory[188] <= 32'h00000000;    //                nop
    memory[189] <= 32'h00000000;    //                nop
    memory[190] <= 32'h00000000;    //                nop
    memory[191] <= 32'h00000000;    //                nop
    memory[192] <= 32'h34047bb0;    //                ori    $a0, $zero, 31664
    memory[193] <= 32'h34057bc0;    //                ori    $a1, $zero, 31680
    memory[194] <= 32'h34067c00;    //                ori    $a2, $zero, 31744
    memory[195] <= 32'h0c00017f;    //                jal    vbsme
    memory[196] <= 32'h00000000;    //                nop
    memory[197] <= 32'h00000000;    //                nop
    memory[198] <= 32'h00000000;    //                nop
    memory[199] <= 32'h00000000;    //                nop
    memory[200] <= 32'h0c00012f;    //                jal    print_result
    memory[201] <= 32'h00000000;    //                nop
    memory[202] <= 32'h00000000;    //                nop
    memory[203] <= 32'h00000000;    //                nop
    memory[204] <= 32'h00000000;    //                nop
    memory[205] <= 32'h34047c40;    //                ori    $a0, $zero, 31808
    memory[206] <= 32'h34057c50;    //                ori    $a1, $zero, 31824
    memory[207] <= 32'h34067c90;    //                ori    $a2, $zero, 31888
    memory[208] <= 32'h0c00017f;    //                jal    vbsme
    memory[209] <= 32'h00000000;    //                nop
    memory[210] <= 32'h00000000;    //                nop
    memory[211] <= 32'h00000000;    //                nop
    memory[212] <= 32'h00000000;    //                nop
    memory[213] <= 32'h0c00012f;    //                jal    print_result
    memory[214] <= 32'h00000000;    //                nop
    memory[215] <= 32'h00000000;    //                nop
    memory[216] <= 32'h00000000;    //                nop
    memory[217] <= 32'h00000000;    //                nop
    memory[218] <= 32'h34047cd8;    //                ori    $a0, $zero, 31960
    memory[219] <= 32'h34057ce8;    //                ori    $a1, $zero, 31976
    memory[220] <= 32'h34067d58;    //                ori    $a2, $zero, 32088
    memory[221] <= 32'h0c00017f;    //                jal    vbsme
    memory[222] <= 32'h00000000;    //                nop
    memory[223] <= 32'h00000000;    //                nop
    memory[224] <= 32'h00000000;    //                nop
    memory[225] <= 32'h00000000;    //                nop
    memory[226] <= 32'h0c00012f;    //                jal    print_result
    memory[227] <= 32'h00000000;    //                nop
    memory[228] <= 32'h00000000;    //                nop
    memory[229] <= 32'h00000000;    //                nop
    memory[230] <= 32'h00000000;    //                nop
    memory[231] <= 32'h34047da0;    //                ori    $a0, $zero, 32160
    memory[232] <= 32'h34057db0;    //                ori    $a1, $zero, 32176
    memory[233] <= 32'h34067e00;    //                ori    $a2, $zero, 32256
    memory[234] <= 32'h0c00017f;    //                jal    vbsme
    memory[235] <= 32'h00000000;    //                nop
    memory[236] <= 32'h00000000;    //                nop
    memory[237] <= 32'h00000000;    //                nop
    memory[238] <= 32'h00000000;    //                nop
    memory[239] <= 32'h0c00012f;    //                jal    print_result
    memory[240] <= 32'h00000000;    //                nop
    memory[241] <= 32'h00000000;    //                nop
    memory[242] <= 32'h00000000;    //                nop
    memory[243] <= 32'h00000000;    //                nop
    memory[244] <= 32'h34047e20;    //                ori    $a0, $zero, 32288
    memory[245] <= 32'h34057e30;    //                ori    $a1, $zero, 32304
    memory[246] <= 32'h34067e80;    //                ori    $a2, $zero, 32384
    memory[247] <= 32'h0c00017f;    //                jal    vbsme
    memory[248] <= 32'h00000000;    //                nop
    memory[249] <= 32'h00000000;    //                nop
    memory[250] <= 32'h00000000;    //                nop
    memory[251] <= 32'h00000000;    //                nop
    memory[252] <= 32'h0c00012f;    //                jal    print_result
    memory[253] <= 32'h00000000;    //                nop
    memory[254] <= 32'h00000000;    //                nop
    memory[255] <= 32'h00000000;    //                nop
    memory[256] <= 32'h00000000;    //                nop
    memory[257] <= 32'h34047e8c;    //                ori    $a0, $zero, 32396
    memory[258] <= 32'h34057e9c;    //                ori    $a1, $zero, 32412
    memory[259] <= 32'h34067eec;    //                ori    $a2, $zero, 32492
    memory[260] <= 32'h0c00017f;    //                jal    vbsme
    memory[261] <= 32'h00000000;    //                nop
    memory[262] <= 32'h00000000;    //                nop
    memory[263] <= 32'h00000000;    //                nop
    memory[264] <= 32'h00000000;    //                nop
    memory[265] <= 32'h0c00012f;    //                jal    print_result
    memory[266] <= 32'h00000000;    //                nop
    memory[267] <= 32'h00000000;    //                nop
    memory[268] <= 32'h00000000;    //                nop
    memory[269] <= 32'h00000000;    //                nop
    memory[270] <= 32'h34047ef8;    //                ori    $a0, $zero, 32504
    memory[271] <= 32'h34057f08;    //                ori    $a1, $zero, 32520
    memory[272] <= 32'h34067f50;    //                ori    $a2, $zero, 32592
    memory[273] <= 32'h0c00017f;    //                jal    vbsme
    memory[274] <= 32'h00000000;    //                nop
    memory[275] <= 32'h00000000;    //                nop
    memory[276] <= 32'h00000000;    //                nop
    memory[277] <= 32'h00000000;    //                nop
    memory[278] <= 32'h0c00012f;    //                jal    print_result
    memory[279] <= 32'h00000000;    //                nop
    memory[280] <= 32'h00000000;    //                nop
    memory[281] <= 32'h00000000;    //                nop
    memory[282] <= 32'h00000000;    //                nop
    memory[283] <= 32'h8fbf0000;    //                lw    $ra, 0($sp)
    memory[284] <= 32'h00000000;    //                nop
    memory[285] <= 32'h00000000;    //                nop
    memory[286] <= 32'h00000000;    //                nop
    memory[287] <= 32'h00000000;    //                nop
    memory[288] <= 32'h23bd0004;    //                addi    $sp, $sp, 4
    memory[289] <= 32'h00000000;    //                nop
    memory[290] <= 32'h00000000;    //                nop
    memory[291] <= 32'h00000000;    //                nop
    memory[292] <= 32'h00000000;    //                nop
    memory[293] <= 32'h3402000a;    //    exit:            ori    $v0, $zero, 10
    memory[294] <= 32'h00000000;    //                nop
    memory[295] <= 32'h00000000;    //                nop
    memory[296] <= 32'h00000000;    //                nop
    memory[297] <= 32'h00000000;    //                nop
    memory[298] <= 32'h00000000;    //                nop
    memory[299] <= 32'h00000000;    //                nop
    memory[300] <= 32'h00000000;    //                nop
    memory[301] <= 32'h00000000;    //                nop
    memory[302] <= 32'h00000000;    //                nop
    memory[303] <= 32'h00402020;    //    print_result:        add    $a0, $v0, $zero
    memory[304] <= 32'h00000000;    //                nop
    memory[305] <= 32'h00000000;    //                nop
    memory[306] <= 32'h00000000;    //                nop
    memory[307] <= 32'h00000000;    //                nop
    memory[308] <= 32'h34020001;    //                ori    $v0, $zero, 1
    memory[309] <= 32'h00000000;    //                nop
    memory[310] <= 32'h00000000;    //                nop
    memory[311] <= 32'h00000000;    //                nop
    memory[312] <= 32'h00000000;    //                nop
    memory[313] <= 32'h00000000;    //                nop
    memory[314] <= 32'h00000000;    //                nop
    memory[315] <= 32'h00000000;    //                nop
    memory[316] <= 32'h00000000;    //                nop
    memory[317] <= 32'h00000000;    //                nop
    memory[318] <= 32'h34047f74;    //                ori    $a0, $zero, 32628
    memory[319] <= 32'h00000000;    //                nop
    memory[320] <= 32'h00000000;    //                nop
    memory[321] <= 32'h00000000;    //                nop
    memory[322] <= 32'h00000000;    //                nop
    memory[323] <= 32'h34020004;    //                ori    $v0, $zero, 4
    memory[324] <= 32'h00000000;    //                nop
    memory[325] <= 32'h00000000;    //                nop
    memory[326] <= 32'h00000000;    //                nop
    memory[327] <= 32'h00000000;    //                nop
    memory[328] <= 32'h00000000;    //                nop
    memory[329] <= 32'h00000000;    //                nop
    memory[330] <= 32'h00000000;    //                nop
    memory[331] <= 32'h00000000;    //                nop
    memory[332] <= 32'h00000000;    //                nop
    memory[333] <= 32'h00602020;    //                add    $a0, $v1, $zero
    memory[334] <= 32'h00000000;    //                nop
    memory[335] <= 32'h00000000;    //                nop
    memory[336] <= 32'h00000000;    //                nop
    memory[337] <= 32'h00000000;    //                nop
    memory[338] <= 32'h34020001;    //                ori    $v0, $zero, 1
    memory[339] <= 32'h00000000;    //                nop
    memory[340] <= 32'h00000000;    //                nop
    memory[341] <= 32'h00000000;    //                nop
    memory[342] <= 32'h00000000;    //                nop
    memory[343] <= 32'h00000000;    //                nop
    memory[344] <= 32'h00000000;    //                nop
    memory[345] <= 32'h00000000;    //                nop
    memory[346] <= 32'h00000000;    //                nop
    memory[347] <= 32'h00000000;    //                nop
    memory[348] <= 32'h34047f74;    //                ori    $a0, $zero, 32628
    memory[349] <= 32'h00000000;    //                nop
    memory[350] <= 32'h00000000;    //                nop
    memory[351] <= 32'h00000000;    //                nop
    memory[352] <= 32'h00000000;    //                nop
    memory[353] <= 32'h34020004;    //                ori    $v0, $zero, 4
    memory[354] <= 32'h00000000;    //                nop
    memory[355] <= 32'h00000000;    //                nop
    memory[356] <= 32'h00000000;    //                nop
    memory[357] <= 32'h00000000;    //                nop
    memory[358] <= 32'h00000000;    //                nop
    memory[359] <= 32'h00000000;    //                nop
    memory[360] <= 32'h00000000;    //                nop
    memory[361] <= 32'h00000000;    //                nop
    memory[362] <= 32'h00000000;    //                nop
    memory[363] <= 32'h34047f74;    //                ori    $a0, $zero, 32628
    memory[364] <= 32'h00000000;    //                nop
    memory[365] <= 32'h00000000;    //                nop
    memory[366] <= 32'h00000000;    //                nop
    memory[367] <= 32'h00000000;    //                nop
    memory[368] <= 32'h34020004;    //                ori    $v0, $zero, 4
    memory[369] <= 32'h00000000;    //                nop
    memory[370] <= 32'h00000000;    //                nop
    memory[371] <= 32'h00000000;    //                nop
    memory[372] <= 32'h00000000;    //                nop
    memory[373] <= 32'h00000000;    //                nop
    memory[374] <= 32'h00000000;    //                nop
    memory[375] <= 32'h00000000;    //                nop
    memory[376] <= 32'h00000000;    //                nop
    memory[377] <= 32'h00000000;    //                nop
    memory[378] <= 32'h03e00008;    //                jr    $ra
    memory[379] <= 32'h00000000;    //                nop
    memory[380] <= 32'h00000000;    //                nop
    memory[381] <= 32'h00000000;    //                nop
    memory[382] <= 32'h00000000;    //                nop
    memory[383] <= 32'h8c900000;    //    vbsme:            lw    $s0, 0($a0)
    memory[384] <= 32'h00000000;    //                nop
    memory[385] <= 32'h00000000;    //                nop
    memory[386] <= 32'h00000000;    //                nop
    memory[387] <= 32'h00000000;    //                nop
    memory[388] <= 32'h8c910004;    //                lw    $s1, 4($a0)
    memory[389] <= 32'h00000000;    //                nop
    memory[390] <= 32'h00000000;    //                nop
    memory[391] <= 32'h00000000;    //                nop
    memory[392] <= 32'h00000000;    //                nop
    memory[393] <= 32'h8c920008;    //                lw    $s2, 8($a0)
    memory[394] <= 32'h00000000;    //                nop
    memory[395] <= 32'h00000000;    //                nop
    memory[396] <= 32'h00000000;    //                nop
    memory[397] <= 32'h00000000;    //                nop
    memory[398] <= 32'h8c93000c;    //                lw    $s3, 12($a0)
    memory[399] <= 32'h00000000;    //                nop
    memory[400] <= 32'h00000000;    //                nop
    memory[401] <= 32'h00000000;    //                nop
    memory[402] <= 32'h00000000;    //                nop
    memory[403] <= 32'h340e0000;    //                ori    $t6, $zero, 0
    memory[404] <= 32'h00000000;    //                nop
    memory[405] <= 32'h00000000;    //                nop
    memory[406] <= 32'h00000000;    //                nop
    memory[407] <= 32'h00000000;    //                nop
    memory[408] <= 32'h340f0000;    //                ori    $t7, $zero, 0
    memory[409] <= 32'h00000000;    //                nop
    memory[410] <= 32'h00000000;    //                nop
    memory[411] <= 32'h00000000;    //                nop
    memory[412] <= 32'h00000000;    //                nop
    memory[413] <= 32'h02124022;    //                sub    $t0, $s0, $s2
    memory[414] <= 32'h00000000;    //                nop
    memory[415] <= 32'h00000000;    //                nop
    memory[416] <= 32'h00000000;    //                nop
    memory[417] <= 32'h00000000;    //                nop
    memory[418] <= 32'h71114002;    //                mul    $t0, $t0, $s1
    memory[419] <= 32'h00000000;    //                nop
    memory[420] <= 32'h00000000;    //                nop
    memory[421] <= 32'h00000000;    //                nop
    memory[422] <= 32'h00000000;    //                nop
    memory[423] <= 32'h02334822;    //                sub    $t1, $s1, $s3
    memory[424] <= 32'h00000000;    //                nop
    memory[425] <= 32'h00000000;    //                nop
    memory[426] <= 32'h00000000;    //                nop
    memory[427] <= 32'h00000000;    //                nop
    memory[428] <= 32'h0109a820;    //                add    $s5, $t0, $t1
    memory[429] <= 32'h00000000;    //                nop
    memory[430] <= 32'h00000000;    //                nop
    memory[431] <= 32'h00000000;    //                nop
    memory[432] <= 32'h00000000;    //                nop
    memory[433] <= 32'hafa80004;    //                sw    $t0, 4($sp)
    memory[434] <= 32'h00000000;    //                nop
    memory[435] <= 32'h00000000;    //                nop
    memory[436] <= 32'h00000000;    //                nop
    memory[437] <= 32'h00000000;    //                nop
    memory[438] <= 32'h34020000;    //                ori    $v0, $zero, 0
    memory[439] <= 32'h00000000;    //                nop
    memory[440] <= 32'h00000000;    //                nop
    memory[441] <= 32'h00000000;    //                nop
    memory[442] <= 32'h00000000;    //                nop
    memory[443] <= 32'h34030000;    //                ori    $v1, $zero, 0
    memory[444] <= 32'h00000000;    //                nop
    memory[445] <= 32'h00000000;    //                nop
    memory[446] <= 32'h00000000;    //                nop
    memory[447] <= 32'h00000000;    //                nop
    memory[448] <= 32'h3416270f;    //                ori    $s6, $zero, 9999
    memory[449] <= 32'h00000000;    //                nop
    memory[450] <= 32'h00000000;    //                nop
    memory[451] <= 32'h00000000;    //                nop
    memory[452] <= 32'h00000000;    //                nop
    memory[453] <= 32'h23bdfffc;    //                addi    $sp, $sp, -4
    memory[454] <= 32'h00000000;    //                nop
    memory[455] <= 32'h00000000;    //                nop
    memory[456] <= 32'h00000000;    //                nop
    memory[457] <= 32'h00000000;    //                nop
    memory[458] <= 32'hafbf0000;    //                sw    $ra, 0($sp)
    memory[459] <= 32'h00000000;    //                nop
    memory[460] <= 32'h00000000;    //                nop
    memory[461] <= 32'h00000000;    //                nop
    memory[462] <= 32'h00000000;    //                nop
    memory[463] <= 32'h0271402a;    //                slt    $t0, $s3, $s1
    memory[464] <= 32'h00000000;    //                nop
    memory[465] <= 32'h00000000;    //                nop
    memory[466] <= 32'h00000000;    //                nop
    memory[467] <= 32'h00000000;    //                nop
    memory[468] <= 32'h0250482a;    //                slt    $t1, $s2, $s0
    memory[469] <= 32'h00000000;    //                nop
    memory[470] <= 32'h00000000;    //                nop
    memory[471] <= 32'h00000000;    //                nop
    memory[472] <= 32'h00000000;    //                nop
    memory[473] <= 32'h01094025;    //                or    $t0, $t0, $t1
    memory[474] <= 32'h00000000;    //                nop
    memory[475] <= 32'h00000000;    //                nop
    memory[476] <= 32'h00000000;    //                nop
    memory[477] <= 32'h00000000;    //                nop
    memory[478] <= 32'h1100012c;    //                beq    $t0, $0, endzigzag
    memory[479] <= 32'h00000000;    //                nop
    memory[480] <= 32'h00000000;    //                nop
    memory[481] <= 32'h00000000;    //                nop
    memory[482] <= 32'h00000000;    //                nop
    memory[483] <= 32'h0c000315;    //                jal    sad
    memory[484] <= 32'h00000000;    //                nop
    memory[485] <= 32'h00000000;    //                nop
    memory[486] <= 32'h00000000;    //                nop
    memory[487] <= 32'h00000000;    //                nop
    memory[488] <= 32'h02334022;    //                sub    $t0, $s1, $s3
    memory[489] <= 32'h00000000;    //                nop
    memory[490] <= 32'h00000000;    //                nop
    memory[491] <= 32'h00000000;    //                nop
    memory[492] <= 32'h00000000;    //                nop
    memory[493] <= 32'h01e8402a;    //                slt    $t0, $t7, $t0
    memory[494] <= 32'h00000000;    //                nop
    memory[495] <= 32'h00000000;    //                nop
    memory[496] <= 32'h00000000;    //                nop
    memory[497] <= 32'h00000000;    //                nop
    memory[498] <= 32'h1100000e;    //                beq    $t0, $0, errordetectnexta
    memory[499] <= 32'h00000000;    //                nop
    memory[500] <= 32'h00000000;    //                nop
    memory[501] <= 32'h00000000;    //                nop
    memory[502] <= 32'h00000000;    //                nop
    memory[503] <= 32'h0c0003c9;    //                jal    rightsubroutine
    memory[504] <= 32'h00000000;    //                nop
    memory[505] <= 32'h00000000;    //                nop
    memory[506] <= 32'h00000000;    //                nop
    memory[507] <= 32'h00000000;    //                nop
    memory[508] <= 32'h08000211;    //                j    doneerrordetectright
    memory[509] <= 32'h00000000;    //                nop
    memory[510] <= 32'h00000000;    //                nop
    memory[511] <= 32'h00000000;    //                nop
    memory[512] <= 32'h00000000;    //                nop
    memory[513] <= 32'h02124022;    //    errordetectnexta:    sub    $t0, $s0, $s2
    memory[514] <= 32'h00000000;    //                nop
    memory[515] <= 32'h00000000;    //                nop
    memory[516] <= 32'h00000000;    //                nop
    memory[517] <= 32'h00000000;    //                nop
    memory[518] <= 32'h01c8402a;    //                slt    $t0, $t6, $t0
    memory[519] <= 32'h00000000;    //                nop
    memory[520] <= 32'h00000000;    //                nop
    memory[521] <= 32'h00000000;    //                nop
    memory[522] <= 32'h00000000;    //                nop
    memory[523] <= 32'h110000ff;    //                beq    $t0, $0, endzigzag
    memory[524] <= 32'h0c0003f1;    //                jal    downsubroutine
    memory[525] <= 32'h00000000;    //                nop
    memory[526] <= 32'h00000000;    //                nop
    memory[527] <= 32'h00000000;    //                nop
    memory[528] <= 32'h00000000;    //                nop
    memory[529] <= 32'h0c000315;    //    doneerrordetectright:    jal    sad
    memory[530] <= 32'h00000000;    //                nop
    memory[531] <= 32'h00000000;    //                nop
    memory[532] <= 32'h00000000;    //                nop
    memory[533] <= 32'h00000000;    //                nop
    memory[534] <= 32'h71d14002;    //    zigzagloop:        mul    $t0, $t6, $s1
    memory[535] <= 32'h00000000;    //                nop
    memory[536] <= 32'h00000000;    //                nop
    memory[537] <= 32'h00000000;    //                nop
    memory[538] <= 32'h00000000;    //                nop
    memory[539] <= 32'h010f4020;    //                add    $t0, $t0, $t7
    memory[540] <= 32'h00000000;    //                nop
    memory[541] <= 32'h00000000;    //                nop
    memory[542] <= 32'h00000000;    //                nop
    memory[543] <= 32'h00000000;    //                nop
    memory[544] <= 32'h0115402a;    //                slt    $t0, $t0, $s5
    memory[545] <= 32'h00000000;    //                nop
    memory[546] <= 32'h00000000;    //                nop
    memory[547] <= 32'h00000000;    //                nop
    memory[548] <= 32'h00000000;    //                nop
    memory[549] <= 32'h110000e5;    //                beq    $t0, $0, endzigzag
    memory[550] <= 32'h00000000;    //                nop
    memory[551] <= 32'h00000000;    //                nop
    memory[552] <= 32'h00000000;    //                nop
    memory[553] <= 32'h00000000;    //                nop
    memory[554] <= 32'h20140001;    //                addi    $s4, $0, 1
    memory[555] <= 32'h00000000;    //                nop
    memory[556] <= 32'h00000000;    //                nop
    memory[557] <= 32'h00000000;    //                nop
    memory[558] <= 32'h00000000;    //                nop
    memory[559] <= 32'h1280004a;    //    dlcollisiondetect:    beq    $s4, $0, edlcollisiondetect
    memory[560] <= 32'h00000000;    //                nop
    memory[561] <= 32'h00000000;    //                nop
    memory[562] <= 32'h00000000;    //                nop
    memory[563] <= 32'h00000000;    //                nop
    memory[564] <= 32'h02124022;    //                sub    $t0, $s0, $s2
    memory[565] <= 32'h00000000;    //                nop
    memory[566] <= 32'h00000000;    //                nop
    memory[567] <= 32'h00000000;    //                nop
    memory[568] <= 32'h00000000;    //                nop
    memory[569] <= 32'h01c8402a;    //                slt    $t0, $t6, $t0
    memory[570] <= 32'h00000000;    //                nop
    memory[571] <= 32'h00000000;    //                nop
    memory[572] <= 32'h00000000;    //                nop
    memory[573] <= 32'h00000000;    //                nop
    memory[574] <= 32'h11000027;    //                beq    $t0, $0, downcollisiona
    memory[575] <= 32'h00000000;    //                nop
    memory[576] <= 32'h00000000;    //                nop
    memory[577] <= 32'h00000000;    //                nop
    memory[578] <= 32'h00000000;    //                nop
    memory[579] <= 32'h000f402a;    //                slt    $t0, $0, $t7
    memory[580] <= 32'h00000000;    //                nop
    memory[581] <= 32'h00000000;    //                nop
    memory[582] <= 32'h00000000;    //                nop
    memory[583] <= 32'h00000000;    //                nop
    memory[584] <= 32'h1100000e;    //                beq    $t0, $0, leftcollisiona
    memory[585] <= 32'h00000000;    //                nop
    memory[586] <= 32'h00000000;    //                nop
    memory[587] <= 32'h00000000;    //                nop
    memory[588] <= 32'h00000000;    //                nop
    memory[589] <= 32'h0c0003d3;    //                jal    downleftsubroutine
    memory[590] <= 32'h00000000;    //                nop
    memory[591] <= 32'h00000000;    //                nop
    memory[592] <= 32'h00000000;    //                nop
    memory[593] <= 32'h00000000;    //                nop
    memory[594] <= 32'h08000270;    //                j    downcollisionaend
    memory[595] <= 32'h00000000;    //                nop
    memory[596] <= 32'h00000000;    //                nop
    memory[597] <= 32'h00000000;    //                nop
    memory[598] <= 32'h00000000;    //                nop
    memory[599] <= 32'h0c0003f1;    //    leftcollisiona:        jal    downsubroutine
    memory[600] <= 32'h00000000;    //                nop
    memory[601] <= 32'h00000000;    //                nop
    memory[602] <= 32'h00000000;    //                nop
    memory[603] <= 32'h00000000;    //                nop
    memory[604] <= 32'h0000a020;    //                add    $s4, $0, $0
    memory[605] <= 32'h00000000;    //                nop
    memory[606] <= 32'h00000000;    //                nop
    memory[607] <= 32'h00000000;    //                nop
    memory[608] <= 32'h00000000;    //                nop
    memory[609] <= 32'h08000270;    //                j    downcollisionaend
    memory[610] <= 32'h00000000;    //                nop
    memory[611] <= 32'h00000000;    //                nop
    memory[612] <= 32'h00000000;    //                nop
    memory[613] <= 32'h00000000;    //                nop
    memory[614] <= 32'h0c0003c9;    //    downcollisiona:        jal    rightsubroutine
    memory[615] <= 32'h00000000;    //                nop
    memory[616] <= 32'h00000000;    //                nop
    memory[617] <= 32'h00000000;    //                nop
    memory[618] <= 32'h00000000;    //                nop
    memory[619] <= 32'h0000a020;    //                add    $s4, $0, $0
    memory[620] <= 32'h00000000;    //                nop
    memory[621] <= 32'h00000000;    //                nop
    memory[622] <= 32'h00000000;    //                nop
    memory[623] <= 32'h00000000;    //                nop
    memory[624] <= 32'h0c000315;    //    downcollisionaend:    jal    sad
    memory[625] <= 32'h00000000;    //                nop
    memory[626] <= 32'h00000000;    //                nop
    memory[627] <= 32'h00000000;    //                nop
    memory[628] <= 32'h00000000;    //                nop
    memory[629] <= 32'h0800022f;    //                j    dlcollisiondetect
    memory[630] <= 32'h00000000;    //                nop
    memory[631] <= 32'h00000000;    //                nop
    memory[632] <= 32'h00000000;    //                nop
    memory[633] <= 32'h00000000;    //                nop
    memory[634] <= 32'h0c000315;    //    edlcollisiondetect:    jal    sad
    memory[635] <= 32'h00000000;    //                nop
    memory[636] <= 32'h00000000;    //                nop
    memory[637] <= 32'h00000000;    //                nop
    memory[638] <= 32'h00000000;    //                nop
    memory[639] <= 32'h71d14002;    //                mul    $t0, $t6, $s1
    memory[640] <= 32'h00000000;    //                nop
    memory[641] <= 32'h00000000;    //                nop
    memory[642] <= 32'h00000000;    //                nop
    memory[643] <= 32'h00000000;    //                nop
    memory[644] <= 32'h010f4020;    //                add    $t0, $t0, $t7
    memory[645] <= 32'h00000000;    //                nop
    memory[646] <= 32'h00000000;    //                nop
    memory[647] <= 32'h00000000;    //                nop
    memory[648] <= 32'h00000000;    //                nop
    memory[649] <= 32'h0115402a;    //                slt    $t0, $t0, $s5
    memory[650] <= 32'h00000000;    //                nop
    memory[651] <= 32'h00000000;    //                nop
    memory[652] <= 32'h00000000;    //                nop
    memory[653] <= 32'h00000000;    //                nop
    memory[654] <= 32'h1100007c;    //                beq    $t0, $0, endzigzag
    memory[655] <= 32'h00000000;    //                nop
    memory[656] <= 32'h00000000;    //                nop
    memory[657] <= 32'h00000000;    //                nop
    memory[658] <= 32'h00000000;    //                nop
    memory[659] <= 32'h20140001;    //                addi    $s4, $0, 1
    memory[660] <= 32'h00000000;    //                nop
    memory[661] <= 32'h00000000;    //                nop
    memory[662] <= 32'h00000000;    //                nop
    memory[663] <= 32'h00000000;    //                nop
    memory[664] <= 32'h12800068;    //    urcollisiondetect:    beq    $s4, $0, eurcollisiondetect
    memory[665] <= 32'h00000000;    //                nop
    memory[666] <= 32'h00000000;    //                nop
    memory[667] <= 32'h00000000;    //                nop
    memory[668] <= 32'h00000000;    //                nop
    memory[669] <= 32'h000e402a;    //                slt    $t0, $0, $t6
    memory[670] <= 32'h00000000;    //                nop
    memory[671] <= 32'h00000000;    //                nop
    memory[672] <= 32'h00000000;    //                nop
    memory[673] <= 32'h00000000;    //                nop
    memory[674] <= 32'h1100002c;    //                beq    $t0, $0, upcollisiona
    memory[675] <= 32'h00000000;    //                nop
    memory[676] <= 32'h00000000;    //                nop
    memory[677] <= 32'h00000000;    //                nop
    memory[678] <= 32'h00000000;    //                nop
    memory[679] <= 32'h02334022;    //                sub    $t0, $s1, $s3
    memory[680] <= 32'h00000000;    //                nop
    memory[681] <= 32'h00000000;    //                nop
    memory[682] <= 32'h00000000;    //                nop
    memory[683] <= 32'h00000000;    //                nop
    memory[684] <= 32'h01e8402a;    //                slt    $t0, $t7, $t0
    memory[685] <= 32'h00000000;    //                nop
    memory[686] <= 32'h00000000;    //                nop
    memory[687] <= 32'h00000000;    //                nop
    memory[688] <= 32'h00000000;    //                nop
    memory[689] <= 32'h1100000e;    //                beq    $t0, $0, rightcollisiona
    memory[690] <= 32'h00000000;    //                nop
    memory[691] <= 32'h00000000;    //                nop
    memory[692] <= 32'h00000000;    //                nop
    memory[693] <= 32'h00000000;    //                nop
    memory[694] <= 32'h0c0003e2;    //                jal    uprightsubroutine
    memory[695] <= 32'h00000000;    //                nop
    memory[696] <= 32'h00000000;    //                nop
    memory[697] <= 32'h00000000;    //                nop
    memory[698] <= 32'h00000000;    //                nop
    memory[699] <= 32'h080002f7;    //                j    upcollisionaend
    memory[700] <= 32'h00000000;    //                nop
    memory[701] <= 32'h00000000;    //                nop
    memory[702] <= 32'h00000000;    //                nop
    memory[703] <= 32'h00000000;    //                nop
    memory[704] <= 32'h0c0003f1;    //    rightcollisiona:    jal    downsubroutine
    memory[705] <= 32'h00000000;    //                nop
    memory[706] <= 32'h00000000;    //                nop
    memory[707] <= 32'h00000000;    //                nop
    memory[708] <= 32'h00000000;    //                nop
    memory[709] <= 32'h0000a020;    //                add    $s4, $0, $0
    memory[710] <= 32'h00000000;    //                nop
    memory[711] <= 32'h00000000;    //                nop
    memory[712] <= 32'h00000000;    //                nop
    memory[713] <= 32'h00000000;    //                nop
    memory[714] <= 32'h080002f7;    //                j    upcollisionaend
    memory[715] <= 32'h00000000;    //                nop
    memory[716] <= 32'h00000000;    //                nop
    memory[717] <= 32'h00000000;    //                nop
    memory[718] <= 32'h00000000;    //                nop
    memory[719] <= 32'h02334022;    //    upcollisiona:        sub    $t0, $s1, $s3
    memory[720] <= 32'h00000000;    //                nop
    memory[721] <= 32'h00000000;    //                nop
    memory[722] <= 32'h00000000;    //                nop
    memory[723] <= 32'h00000000;    //                nop
    memory[724] <= 32'h01e8402a;    //                slt    $t0, $t7, $t0
    memory[725] <= 32'h00000000;    //                nop
    memory[726] <= 32'h00000000;    //                nop
    memory[727] <= 32'h00000000;    //                nop
    memory[728] <= 32'h00000000;    //                nop
    memory[729] <= 32'h11000013;    //                beq    $t0, $0, rightcollisionb
    memory[730] <= 32'h00000000;    //                nop
    memory[731] <= 32'h00000000;    //                nop
    memory[732] <= 32'h00000000;    //                nop
    memory[733] <= 32'h00000000;    //                nop
    memory[734] <= 32'h0c0003c9;    //                jal    rightsubroutine
    memory[735] <= 32'h00000000;    //                nop
    memory[736] <= 32'h00000000;    //                nop
    memory[737] <= 32'h00000000;    //                nop
    memory[738] <= 32'h00000000;    //                nop
    memory[739] <= 32'h0000a020;    //                add    $s4, $0, $0
    memory[740] <= 32'h00000000;    //                nop
    memory[741] <= 32'h00000000;    //                nop
    memory[742] <= 32'h00000000;    //                nop
    memory[743] <= 32'h00000000;    //                nop
    memory[744] <= 32'h080002f7;    //                j    upcollisionaend
    memory[745] <= 32'h00000000;    //                nop
    memory[746] <= 32'h00000000;    //                nop
    memory[747] <= 32'h00000000;    //                nop
    memory[748] <= 32'h00000000;    //                nop
    memory[749] <= 32'h0c0003f1;    //    rightcollisionb:    jal    downsubroutine
    memory[750] <= 32'h00000000;    //                nop
    memory[751] <= 32'h00000000;    //                nop
    memory[752] <= 32'h00000000;    //                nop
    memory[753] <= 32'h00000000;    //                nop
    memory[754] <= 32'h0000a020;    //                add    $s4, $0, $0
    memory[755] <= 32'h00000000;    //                nop
    memory[756] <= 32'h00000000;    //                nop
    memory[757] <= 32'h00000000;    //                nop
    memory[758] <= 32'h00000000;    //                nop
    memory[759] <= 32'h0c000315;    //    upcollisionaend:    jal    sad
    memory[760] <= 32'h00000000;    //                nop
    memory[761] <= 32'h00000000;    //                nop
    memory[762] <= 32'h00000000;    //                nop
    memory[763] <= 32'h00000000;    //                nop
    memory[764] <= 32'h08000298;    //                j    urcollisiondetect
    memory[765] <= 32'h00000000;    //                nop
    memory[766] <= 32'h00000000;    //                nop
    memory[767] <= 32'h00000000;    //                nop
    memory[768] <= 32'h00000000;    //                nop
    memory[769] <= 32'h0c000315;    //    eurcollisiondetect:    jal    sad
    memory[770] <= 32'h00000000;    //                nop
    memory[771] <= 32'h00000000;    //                nop
    memory[772] <= 32'h00000000;    //                nop
    memory[773] <= 32'h00000000;    //                nop
    memory[774] <= 32'h08000216;    //                j    zigzagloop
    memory[775] <= 32'h00000000;    //                nop
    memory[776] <= 32'h00000000;    //                nop
    memory[777] <= 32'h00000000;    //                nop
    memory[778] <= 32'h00000000;    //                nop
    memory[779] <= 32'h8fbf0000;    //    endzigzag:        lw    $ra, 0($sp)
    memory[780] <= 32'h00000000;    //                nop
    memory[781] <= 32'h00000000;    //                nop
    memory[782] <= 32'h00000000;    //                nop
    memory[783] <= 32'h00000000;    //                nop
    memory[784] <= 32'h03e00008;    //                jr    $ra
    memory[785] <= 32'h00000000;    //                nop
    memory[786] <= 32'h00000000;    //                nop
    memory[787] <= 32'h00000000;    //                nop
    memory[788] <= 32'h00000000;    //                nop
    memory[789] <= 32'h00004020;    //    sad:            add    $t0, $0, $0
    memory[790] <= 32'h00000000;    //                nop
    memory[791] <= 32'h00000000;    //                nop
    memory[792] <= 32'h00000000;    //                nop
    memory[793] <= 32'h00000000;    //                nop
    memory[794] <= 32'h00004820;    //                add    $t1, $0, $0
    memory[795] <= 32'h00000000;    //                nop
    memory[796] <= 32'h00000000;    //                nop
    memory[797] <= 32'h00000000;    //                nop
    memory[798] <= 32'h00000000;    //                nop
    memory[799] <= 32'h0132582a;    //    sadouterloop:        slt    $t3, $t1, $s2
    memory[800] <= 32'h00000000;    //                nop
    memory[801] <= 32'h00000000;    //                nop
    memory[802] <= 32'h00000000;    //                nop
    memory[803] <= 32'h00000000;    //                nop
    memory[804] <= 32'h11600081;    //                beq    $t3, $0, sadouterloopend
    memory[805] <= 32'h00000000;    //                nop
    memory[806] <= 32'h00000000;    //                nop
    memory[807] <= 32'h00000000;    //                nop
    memory[808] <= 32'h00000000;    //                nop
    memory[809] <= 32'h00005020;    //                add    $t2, $0, $0
    memory[810] <= 32'h00000000;    //                nop
    memory[811] <= 32'h00000000;    //                nop
    memory[812] <= 32'h00000000;    //                nop
    memory[813] <= 32'h00000000;    //                nop
    memory[814] <= 32'h0153582a;    //    sadinnerloop:        slt    $t3, $t2, $s3
    memory[815] <= 32'h00000000;    //                nop
    memory[816] <= 32'h00000000;    //                nop
    memory[817] <= 32'h00000000;    //                nop
    memory[818] <= 32'h00000000;    //                nop
    memory[819] <= 32'h11600068;    //                beq    $t3, $0, sadinnerloopend
    memory[820] <= 32'h00000000;    //                nop
    memory[821] <= 32'h00000000;    //                nop
    memory[822] <= 32'h00000000;    //                nop
    memory[823] <= 32'h00000000;    //                nop
    memory[824] <= 32'h012e5820;    //                add    $t3, $t1, $t6
    memory[825] <= 32'h00000000;    //                nop
    memory[826] <= 32'h00000000;    //                nop
    memory[827] <= 32'h00000000;    //                nop
    memory[828] <= 32'h00000000;    //                nop
    memory[829] <= 32'h71715802;    //                mul    $t3, $t3, $s1
    memory[830] <= 32'h00000000;    //                nop
    memory[831] <= 32'h00000000;    //                nop
    memory[832] <= 32'h00000000;    //                nop
    memory[833] <= 32'h00000000;    //                nop
    memory[834] <= 32'h016a5820;    //                add    $t3, $t3, $t2
    memory[835] <= 32'h00000000;    //                nop
    memory[836] <= 32'h00000000;    //                nop
    memory[837] <= 32'h00000000;    //                nop
    memory[838] <= 32'h00000000;    //                nop
    memory[839] <= 32'h016f5820;    //                add    $t3, $t3, $t7
    memory[840] <= 32'h00000000;    //                nop
    memory[841] <= 32'h00000000;    //                nop
    memory[842] <= 32'h00000000;    //                nop
    memory[843] <= 32'h00000000;    //                nop
    memory[844] <= 32'h000b5880;    //                sll    $t3, $t3, 2
    memory[845] <= 32'h00000000;    //                nop
    memory[846] <= 32'h00000000;    //                nop
    memory[847] <= 32'h00000000;    //                nop
    memory[848] <= 32'h00000000;    //                nop
    memory[849] <= 32'h71336002;    //                mul    $t4, $t1, $s3
    memory[850] <= 32'h00000000;    //                nop
    memory[851] <= 32'h00000000;    //                nop
    memory[852] <= 32'h00000000;    //                nop
    memory[853] <= 32'h00000000;    //                nop
    memory[854] <= 32'h018a6020;    //                add    $t4, $t4, $t2
    memory[855] <= 32'h00000000;    //                nop
    memory[856] <= 32'h00000000;    //                nop
    memory[857] <= 32'h00000000;    //                nop
    memory[858] <= 32'h00000000;    //                nop
    memory[859] <= 32'h000c6080;    //                sll    $t4, $t4, 2
    memory[860] <= 32'h00000000;    //                nop
    memory[861] <= 32'h00000000;    //                nop
    memory[862] <= 32'h00000000;    //                nop
    memory[863] <= 32'h00000000;    //                nop
    memory[864] <= 32'h00ab5820;    //                add    $t3, $a1, $t3
    memory[865] <= 32'h00000000;    //                nop
    memory[866] <= 32'h00000000;    //                nop
    memory[867] <= 32'h00000000;    //                nop
    memory[868] <= 32'h00000000;    //                nop
    memory[869] <= 32'h00cc6020;    //                add    $t4, $a2, $t4
    memory[870] <= 32'h00000000;    //                nop
    memory[871] <= 32'h00000000;    //                nop
    memory[872] <= 32'h00000000;    //                nop
    memory[873] <= 32'h00000000;    //                nop
    memory[874] <= 32'h8d6b0000;    //                lw    $t3, 0($t3)
    memory[875] <= 32'h00000000;    //                nop
    memory[876] <= 32'h00000000;    //                nop
    memory[877] <= 32'h00000000;    //                nop
    memory[878] <= 32'h00000000;    //                nop
    memory[879] <= 32'h8d8c0000;    //                lw    $t4, 0($t4)
    memory[880] <= 32'h00000000;    //                nop
    memory[881] <= 32'h00000000;    //                nop
    memory[882] <= 32'h00000000;    //                nop
    memory[883] <= 32'h00000000;    //                nop
    memory[884] <= 32'h016c5822;    //                sub    $t3, $t3, $t4
    memory[885] <= 32'h00000000;    //                nop
    memory[886] <= 32'h00000000;    //                nop
    memory[887] <= 32'h00000000;    //                nop
    memory[888] <= 32'h00000000;    //                nop
    memory[889] <= 32'h0160602a;    //                slt    $t4, $t3, $0
    memory[890] <= 32'h00000000;    //                nop
    memory[891] <= 32'h00000000;    //                nop
    memory[892] <= 32'h00000000;    //                nop
    memory[893] <= 32'h00000000;    //                nop
    memory[894] <= 32'h1180000e;    //                beq    $t4, $0, absifend
    memory[895] <= 32'h00000000;    //                nop
    memory[896] <= 32'h00000000;    //                nop
    memory[897] <= 32'h00000000;    //                nop
    memory[898] <= 32'h00000000;    //                nop
    memory[899] <= 32'h200dffff;    //                addi    $t5, $0, -1
    memory[900] <= 32'h00000000;    //                nop
    memory[901] <= 32'h00000000;    //                nop
    memory[902] <= 32'h00000000;    //                nop
    memory[903] <= 32'h00000000;    //                nop
    memory[904] <= 32'h716d5802;    //                mul    $t3, $t3, $t5
    memory[905] <= 32'h00000000;    //                nop
    memory[906] <= 32'h00000000;    //                nop
    memory[907] <= 32'h00000000;    //                nop
    memory[908] <= 32'h00000000;    //                nop
    memory[909] <= 32'h010b4020;    //    absifend:        add    $t0, $t0, $t3
    memory[910] <= 32'h00000000;    //                nop
    memory[911] <= 32'h00000000;    //                nop
    memory[912] <= 32'h00000000;    //                nop
    memory[913] <= 32'h00000000;    //                nop
    memory[914] <= 32'h214a0001;    //                addi    $t2, $t2, 1
    memory[915] <= 32'h00000000;    //                nop
    memory[916] <= 32'h00000000;    //                nop
    memory[917] <= 32'h00000000;    //                nop
    memory[918] <= 32'h00000000;    //                nop
    memory[919] <= 32'h0800032e;    //                j    sadinnerloop
    memory[920] <= 32'h00000000;    //                nop
    memory[921] <= 32'h00000000;    //                nop
    memory[922] <= 32'h00000000;    //                nop
    memory[923] <= 32'h00000000;    //                nop
    memory[924] <= 32'h21290001;    //    sadinnerloopend:    addi    $t1, $t1, 1
    memory[925] <= 32'h00000000;    //                nop
    memory[926] <= 32'h00000000;    //                nop
    memory[927] <= 32'h00000000;    //                nop
    memory[928] <= 32'h00000000;    //                nop
    memory[929] <= 32'h0800031f;    //                j    sadouterloop
    memory[930] <= 32'h00000000;    //                nop
    memory[931] <= 32'h00000000;    //                nop
    memory[932] <= 32'h00000000;    //                nop
    memory[933] <= 32'h00000000;    //                nop
    memory[934] <= 32'h1116000e;    //    sadouterloopend:    beq    $t0, $s6, lteqcurrmin
    memory[935] <= 32'h00000000;    //                nop
    memory[936] <= 32'h00000000;    //                nop
    memory[937] <= 32'h00000000;    //                nop
    memory[938] <= 32'h00000000;    //                nop
    memory[939] <= 32'h0116482a;    //                slt    $t1, $t0, $s6
    memory[940] <= 32'h00000000;    //                nop
    memory[941] <= 32'h00000000;    //                nop
    memory[942] <= 32'h00000000;    //                nop
    memory[943] <= 32'h00000000;    //                nop
    memory[944] <= 32'h11200013;    //                beq    $t1, $0, lteqcurrminend
    memory[945] <= 32'h00000000;    //                nop
    memory[946] <= 32'h00000000;    //                nop
    memory[947] <= 32'h00000000;    //                nop
    memory[948] <= 32'h00000000;    //                nop
    memory[949] <= 32'h0100b020;    //    lteqcurrmin:        add    $s6, $t0, $0
    memory[950] <= 32'h00000000;    //                nop
    memory[951] <= 32'h00000000;    //                nop
    memory[952] <= 32'h00000000;    //                nop
    memory[953] <= 32'h00000000;    //                nop
    memory[954] <= 32'h01c01020;    //                add    $v0, $t6, $0
    memory[955] <= 32'h00000000;    //                nop
    memory[956] <= 32'h00000000;    //                nop
    memory[957] <= 32'h00000000;    //                nop
    memory[958] <= 32'h00000000;    //                nop
    memory[959] <= 32'h01e01820;    //                add    $v1, $t7, $0
    memory[960] <= 32'h00000000;    //                nop
    memory[961] <= 32'h00000000;    //                nop
    memory[962] <= 32'h00000000;    //                nop
    memory[963] <= 32'h00000000;    //                nop
    memory[964] <= 32'h03e00008;    //    lteqcurrminend:        jr    $ra
    memory[965] <= 32'h00000000;    //                nop
    memory[966] <= 32'h00000000;    //                nop
    memory[967] <= 32'h00000000;    //                nop
    memory[968] <= 32'h00000000;    //                nop
    memory[969] <= 32'h21ef0001;    //    rightsubroutine:    addi    $t7, $t7, 1
    memory[970] <= 32'h00000000;    //                nop
    memory[971] <= 32'h00000000;    //                nop
    memory[972] <= 32'h00000000;    //                nop
    memory[973] <= 32'h00000000;    //                nop
    memory[974] <= 32'h03e00008;    //                jr    $ra
    memory[975] <= 32'h00000000;    //                nop
    memory[976] <= 32'h00000000;    //                nop
    memory[977] <= 32'h00000000;    //                nop
    memory[978] <= 32'h00000000;    //                nop
    memory[979] <= 32'h21ce0001;    //    downleftsubroutine:    addi    $t6, $t6, 1
    memory[980] <= 32'h00000000;    //                nop
    memory[981] <= 32'h00000000;    //                nop
    memory[982] <= 32'h00000000;    //                nop
    memory[983] <= 32'h00000000;    //                nop
    memory[984] <= 32'h21efffff;    //                addi    $t7, $t7, -1
    memory[985] <= 32'h00000000;    //                nop
    memory[986] <= 32'h00000000;    //                nop
    memory[987] <= 32'h00000000;    //                nop
    memory[988] <= 32'h00000000;    //                nop
    memory[989] <= 32'h03e00008;    //                jr    $ra
    memory[990] <= 32'h00000000;    //                nop
    memory[991] <= 32'h00000000;    //                nop
    memory[992] <= 32'h00000000;    //                nop
    memory[993] <= 32'h00000000;    //                nop
    memory[994] <= 32'h21ceffff;    //    uprightsubroutine:    addi    $t6, $t6, -1
    memory[995] <= 32'h00000000;    //                nop
    memory[996] <= 32'h00000000;    //                nop
    memory[997] <= 32'h00000000;    //                nop
    memory[998] <= 32'h00000000;    //                nop
    memory[999] <= 32'h21ef0001;    //                addi    $t7, $t7, 1
    memory[1000] <= 32'h00000000;    //                nop
    memory[1001] <= 32'h00000000;    //                nop
    memory[1002] <= 32'h00000000;    //                nop
    memory[1003] <= 32'h00000000;    //                nop
    memory[1004] <= 32'h03e00008;    //                jr    $ra
    memory[1005] <= 32'h00000000;    //                nop
    memory[1006] <= 32'h00000000;    //                nop
    memory[1007] <= 32'h00000000;    //                nop
    memory[1008] <= 32'h00000000;    //                nop
    memory[1009] <= 32'h21ce0001;    //    downsubroutine:        addi    $t6, $t6, 1
    memory[1010] <= 32'h00000000;    //                nop
    memory[1011] <= 32'h00000000;    //                nop
    memory[1012] <= 32'h00000000;    //                nop
    memory[1013] <= 32'h00000000;    //                nop
    memory[1014] <= 32'h03e00008;    //                jr    $ra
    memory[1015] <= 32'h00000000;    //                nop
    memory[1016] <= 32'h00000000;    //                nop
    memory[1017] <= 32'h00000000;    //                nop
    memory[1018] <= 32'h00000000;    //                nop
    memory[1019] <= 32'h21ceffff;    //    upsubroutine:        addi    $t6, $t6, -1
    memory[1020] <= 32'h00000000;    //                nop
    memory[1021] <= 32'h00000000;    //                nop
    memory[1022] <= 32'h00000000;    //                nop
    memory[1023] <= 32'h21ef0001;    //                addi    $t7, $t7, 1
    
    */
    
    
    
    
    
    
    
    
    

////        The intermet
//    Memory[0] = 32'h20090006;	//		addi	$t1, $zero, 6
//	Memory[1] = 32'h00000000;	//		nop
//	Memory[2] = 32'h00000000;	//		nop
//	Memory[3] = 32'h00000000;	//		nop
//	Memory[4] = 32'h00000000;	//		nop
//	Memory[5] = 32'h00000000;	//		nop
//	Memory[6] = 32'h200a0008;	//		addi	$t2, $zero, 8
//	Memory[7] = 32'h00000000;	//		nop
//	Memory[8] = 32'h00000000;	//		nop
//	Memory[9] = 32'h00000000;	//		nop
//	Memory[10] = 32'h00000000;	//		nop
//	Memory[11] = 32'h00000000;	//		nop
//	Memory[12] = 32'h01495822;	//		sub	$t3, $t2, $t1
//	Memory[13] = 32'h00000000;	//		nop
//	Memory[14] = 32'h00000000;	//		nop
//	Memory[15] = 32'h00000000;	//		nop
//	Memory[16] = 32'h00000000;	//		nop
//	Memory[17] = 32'h00000000;	//		nop
//	Memory[18] = 32'h000b60c0;	//		sll	$t4, $t3, 3
//	Memory[19] = 32'h00000000;	//		nop
//	Memory[20] = 32'h00000000;	//		nop
//	Memory[21] = 32'h00000000;	//		nop
//	Memory[22] = 32'h00000000;	//		nop
//	Memory[23] = 32'h00000000;	//		nop
//	Memory[24] = 32'h000c6882;	//		srl	$t5, $t4, 2


            

            












/*
//Public Test Case Labs 15-18
memory[0] <= 32'h34040000;	//	        main:		ori	$a0, $zero, 0
memory[1] <= 32'h00000000;	//			nop
memory[2] <= 32'h00000000;	//			nop
memory[3] <= 32'h00000000;	//			nop
memory[4] <= 32'h00000000;	//			nop
memory[5] <= 32'h00000000;	//			nop
memory[6] <= 32'h08000018;	//			j	start
memory[7] <= 32'h00000000;	//			nop
memory[8] <= 32'h00000000;	//			nop
memory[9] <= 32'h00000000;	//			nop
memory[10] <= 32'h00000000;	//			nop
memory[11] <= 32'h00000000;	//			nop
memory[12] <= 32'h2004000a;	//			addi	$a0, $zero, 10
memory[13] <= 32'h00000000;	//			nop
memory[14] <= 32'h00000000;	//			nop
memory[15] <= 32'h00000000;	//			nop
memory[16] <= 32'h00000000;	//			nop
memory[17] <= 32'h00000000;	//			nop
memory[18] <= 32'h2004000a;	//			addi	$a0, $zero, 10
memory[19] <= 32'h00000000;	//			nop
memory[20] <= 32'h00000000;	//			nop
memory[21] <= 32'h00000000;	//			nop
memory[22] <= 32'h00000000;	//			nop
memory[23] <= 32'h00000000;	//			nop
memory[24] <= 32'h8c900004;	//	start:		lw	$s0, 4($a0)
memory[25] <= 32'h00000000;	//			nop        
memory[26] <= 32'h00000000;	//			nop
memory[27] <= 32'h00000000;	//			nop
memory[28] <= 32'h00000000;	//			nop
memory[29] <= 32'h00000000;	//			nop
memory[30] <= 32'h8c900008;	//			lw	$s0, 8($a0)
memory[31] <= 32'h00000000;	//			nop  
memory[32] <= 32'h00000000;	//			nop
memory[33] <= 32'h00000000;	//			nop
memory[34] <= 32'h00000000;	//			nop
memory[35] <= 32'h00000000;	//			nop
memory[36] <= 32'hac900000;	//			sw	$s0, 0($a0)
memory[37] <= 32'h00000000;	//			nop
memory[38] <= 32'h00000000;	//			nop
memory[39] <= 32'h00000000;	//			nop
memory[40] <= 32'h00000000;	//			nop
memory[41] <= 32'h00000000;	//			nop
memory[42] <= 32'hac90000c;	//			sw	$s0, 12($a0)
memory[43] <= 32'h00000000;	//			nop
memory[44] <= 32'h00000000;	//			nop
memory[45] <= 32'h00000000;	//			nop
memory[46] <= 32'h00000000;	//			nop
memory[47] <= 32'h00000000;	//			nop
memory[48] <= 32'h8c910000;	//			lw	$s1, 0($a0)
memory[49] <= 32'h00000000;	//			nop
memory[50] <= 32'h00000000;	//			nop
memory[51] <= 32'h00000000;	//			nop
memory[52] <= 32'h00000000;	//			nop
memory[53] <= 32'h00000000;	//			nop
memory[54] <= 32'h8c92000c;	//			lw	$s2, 12($a0)
memory[55] <= 32'h00000000;	//			nop
memory[56] <= 32'h00000000;	//			nop
memory[57] <= 32'h00000000;	//			nop
memory[58] <= 32'h00000000;	//			nop
memory[59] <= 32'h00000000;	//			nop
memory[60] <= 32'h12000017;	//			beq	$s0, $zero, branch1
memory[61] <= 32'h00000000;	//			nop
memory[62] <= 32'h00000000;	//			nop
memory[63] <= 32'h00000000;	//			nop
memory[64] <= 32'h00000000;	//			nop
memory[65] <= 32'h00000000;	//			nop
memory[66] <= 32'h02008820;	//			add	$s1, $s0, $zero
memory[67] <= 32'h00000000;	//			nop
memory[68] <= 32'h00000000;	//			nop
memory[69] <= 32'h00000000;	//			nop
memory[70] <= 32'h00000000;	//			nop
memory[71] <= 32'h00000000;	//			nop
memory[72] <= 32'h1211000b;	//			beq	$s0, $s1, branch1
memory[73] <= 32'h00000000;	//			nop
memory[74] <= 32'h00000000;	//			nop
memory[75] <= 32'h00000000;	//			nop
memory[76] <= 32'h00000000;	//			nop
memory[77] <= 32'h00000000;	//			nop
memory[78] <= 32'h0800013e;	//			j	error
memory[79] <= 32'h00000000;	//			nop
memory[80] <= 32'h00000000;	//			nop
memory[81] <= 32'h00000000;	//			nop
memory[82] <= 32'h00000000;	//			nop
memory[83] <= 32'h00000000;	//			nop
memory[84] <= 32'h2010ffff;	//	branch1:	addi	$s0, $zero, -1
memory[85] <= 32'h00000000;	//			nop
memory[86] <= 32'h00000000;	//			nop
memory[87] <= 32'h00000000;	//			nop
memory[88] <= 32'h00000000;	//			nop
memory[89] <= 32'h00000000;	//			nop
memory[90] <= 32'h0601ffbd;	//			bgez	$s0, start
memory[91] <= 32'h00000000;	//			nop
memory[92] <= 32'h00000000;	//			nop
memory[93] <= 32'h00000000;	//			nop
memory[94] <= 32'h00000000;	//			nop
memory[95] <= 32'h00000000;	//			nop
memory[96] <= 32'h22100001;	//			addi	$s0, $s0, 1
memory[97] <= 32'h00000000;	//			nop
memory[98] <= 32'h00000000;	//			nop
memory[99] <= 32'h00000000;	//			nop
memory[100] <= 32'h00000000;	//			nop
memory[101] <= 32'h00000000;	//			nop
memory[102] <= 32'h0601000b;	//			bgez	$s0, branch2
memory[103] <= 32'h00000000;	//			nop
memory[104] <= 32'h00000000;	//			nop
memory[105] <= 32'h00000000;	//			nop
memory[106] <= 32'h00000000;	//			nop
memory[107] <= 32'h00000000;	//			nop
memory[108] <= 32'h0800013e;	//			j	error
memory[109] <= 32'h00000000;	//			nop
memory[110] <= 32'h00000000;	//			nop
memory[111] <= 32'h00000000;	//			nop
memory[112] <= 32'h00000000;	//			nop
memory[113] <= 32'h00000000;	//			nop
memory[114] <= 32'h2010ffff;	//	branch2:	addi	$s0, $zero, -1
memory[115] <= 32'h00000000;	//			nop
memory[116] <= 32'h00000000;	//			nop
memory[117] <= 32'h00000000;	//			nop
memory[118] <= 32'h00000000;	//			nop
memory[119] <= 32'h00000000;	//			nop
memory[120] <= 32'h1e000017;	//			bgtz	$s0, branch3
memory[121] <= 32'h00000000;	//			nop
memory[122] <= 32'h00000000;	//			nop
memory[123] <= 32'h00000000;	//			nop
memory[124] <= 32'h00000000;	//			nop
memory[125] <= 32'h00000000;	//			nop
memory[126] <= 32'h20100001;	//			addi	$s0, $zero, 1
memory[127] <= 32'h00000000;	//			nop
memory[128] <= 32'h00000000;	//			nop
memory[129] <= 32'h00000000;	//			nop
memory[130] <= 32'h00000000;	//			nop
memory[131] <= 32'h00000000;	//			nop
memory[132] <= 32'h1e00000b;	//			bgtz	$s0, branch3
memory[133] <= 32'h00000000;	//			nop
memory[134] <= 32'h00000000;	//			nop
memory[135] <= 32'h00000000;	//			nop
memory[136] <= 32'h00000000;	//			nop
memory[137] <= 32'h00000000;	//			nop
memory[138] <= 32'h0800013e;	//			j	error
memory[139] <= 32'h00000000;	//			nop
memory[140] <= 32'h00000000;	//			nop
memory[141] <= 32'h00000000;	//			nop
memory[142] <= 32'h00000000;	//			nop
memory[143] <= 32'h00000000;	//			nop
memory[144] <= 32'h06000017;	//	branch3:	bltz	$s0, branch4
memory[145] <= 32'h00000000;	//			nop
memory[146] <= 32'h00000000;	//			nop
memory[147] <= 32'h00000000;	//			nop
memory[148] <= 32'h00000000;	//			nop
memory[149] <= 32'h00000000;	//			nop
memory[150] <= 32'h2010ffff;	//			addi	$s0, $zero, -1
memory[151] <= 32'h00000000;	//			nop
memory[152] <= 32'h00000000;	//			nop
memory[153] <= 32'h00000000;	//			nop
memory[154] <= 32'h00000000;	//			nop
memory[155] <= 32'h00000000;	//			nop
memory[156] <= 32'h0600000b;	//			bltz	$s0, branch4
memory[157] <= 32'h00000000;	//			nop
memory[158] <= 32'h00000000;	//			nop
memory[159] <= 32'h00000000;	//			nop
memory[160] <= 32'h00000000;	//			nop
memory[161] <= 32'h00000000;	//			nop
memory[162] <= 32'h0800013e;	//			j	error
memory[163] <= 32'h00000000;	//			nop
memory[164] <= 32'h00000000;	//			nop
memory[165] <= 32'h00000000;	//			nop
memory[166] <= 32'h00000000;	//			nop
memory[167] <= 32'h00000000;	//			nop
memory[168] <= 32'h2011ffff;	//	branch4:	addi	$s1, $zero, -1
memory[169] <= 32'h00000000;	//			nop
memory[170] <= 32'h00000000;	//			nop
memory[171] <= 32'h00000000;	//			nop
memory[172] <= 32'h00000000;	//			nop
memory[173] <= 32'h00000000;	//			nop
memory[174] <= 32'h16110011;	//			bne	$s0, $s1, branch5
memory[175] <= 32'h00000000;	//			nop
memory[176] <= 32'h00000000;	//			nop
memory[177] <= 32'h00000000;	//			nop
memory[178] <= 32'h00000000;	//			nop
memory[179] <= 32'h00000000;	//			nop
memory[180] <= 32'h1600000b;	//			bne	$s0, $zero, branch5
memory[181] <= 32'h00000000;	//			nop
memory[182] <= 32'h00000000;	//			nop
memory[183] <= 32'h00000000;	//			nop
memory[184] <= 32'h00000000;	//			nop
memory[185] <= 32'h00000000;	//			nop
memory[186] <= 32'h0800013e;	//			j	error
memory[187] <= 32'h00000000;	//			nop
memory[188] <= 32'h00000000;	//			nop
memory[189] <= 32'h00000000;	//			nop
memory[190] <= 32'h00000000;	//			nop
memory[191] <= 32'h00000000;	//			nop
memory[192] <= 32'h20100080;	//	branch5:	addi	$s0, $zero, 128
memory[193] <= 32'h00000000;	//			nop
memory[194] <= 32'h00000000;	//			nop
memory[195] <= 32'h00000000;	//			nop
memory[196] <= 32'h00000000;	//			nop
memory[197] <= 32'h00000000;	//			nop
memory[198] <= 32'ha0900000;	//			sb	$s0, 0($a0)
memory[199] <= 32'h00000000;	//			nop
memory[200] <= 32'h00000000;	//			nop
memory[201] <= 32'h00000000;	//			nop
memory[202] <= 32'h00000000;	//			nop
memory[203] <= 32'h00000000;	//			nop
memory[204] <= 32'h80900000;	//			lb	$s0, 0($a0)
memory[205] <= 32'h00000000;	//			nop
memory[206] <= 32'h00000000;	//			nop
memory[207] <= 32'h00000000;	//			nop
memory[208] <= 32'h00000000;	//			nop
memory[209] <= 32'h00000000;	//			nop
memory[210] <= 32'h1a00000b;	//			blez	$s0, branch6
memory[211] <= 32'h00000000;	//			nop
memory[212] <= 32'h00000000;	//			nop
memory[213] <= 32'h00000000;	//			nop
memory[214] <= 32'h00000000;	//			nop
memory[215] <= 32'h00000000;	//			nop
memory[216] <= 32'h0800013e;	//			j	error
memory[217] <= 32'h00000000;	//			nop
memory[218] <= 32'h00000000;	//			nop
memory[219] <= 32'h00000000;	//			nop
memory[220] <= 32'h00000000;	//			nop
memory[221] <= 32'h00000000;	//			nop
memory[222] <= 32'h2010ffff;	//	branch6:	addi	$s0, $zero, -1
memory[223] <= 32'h00000000;	//			nop
memory[224] <= 32'h00000000;	//			nop
memory[225] <= 32'h00000000;	//			nop
memory[226] <= 32'h00000000;	//			nop
memory[227] <= 32'h00000000;	//			nop
memory[228] <= 32'ha4900000;	//			sh	$s0, 0($a0)
memory[229] <= 32'h00000000;	//			nop
memory[230] <= 32'h00000000;	//			nop
memory[231] <= 32'h00000000;	//			nop
memory[232] <= 32'h00000000;	//			nop
memory[233] <= 32'h00000000;	//			nop
memory[234] <= 32'h20100000;	//			addi	$s0, $zero, 0
memory[235] <= 32'h00000000;	//			nop
memory[236] <= 32'h00000000;	//			nop
memory[237] <= 32'h00000000;	//			nop
memory[238] <= 32'h00000000;	//			nop
memory[239] <= 32'h00000000;	//			nop
memory[240] <= 32'h84900000;	//			lh	$s0, 0($a0)
memory[241] <= 32'h00000000;	//			nop
memory[242] <= 32'h00000000;	//			nop
memory[243] <= 32'h00000000;	//			nop
memory[244] <= 32'h00000000;	//			nop
memory[245] <= 32'h00000000;	//			nop
memory[246] <= 32'h1a00000b;	//			blez	$s0, branch7
memory[247] <= 32'h00000000;	//			nop
memory[248] <= 32'h00000000;	//			nop
memory[249] <= 32'h00000000;	//			nop
memory[250] <= 32'h00000000;	//			nop
memory[251] <= 32'h00000000;	//			nop
memory[252] <= 32'h0800013e;	//			j	error
memory[253] <= 32'h00000000;	//			nop
memory[254] <= 32'h00000000;	//			nop
memory[255] <= 32'h00000000;	//			nop
memory[256] <= 32'h00000000;	//			nop
memory[257] <= 32'h00000000;	//			nop
memory[258] <= 32'h2010ffff;	//	branch7:	addi	$s0, $zero, -1
memory[259] <= 32'h00000000;	//			nop
memory[260] <= 32'h00000000;	//			nop
memory[261] <= 32'h00000000;	//			nop
memory[262] <= 32'h00000000;	//			nop
memory[263] <= 32'h00000000;	//			nop
memory[264] <= 32'h3c100001;	//			lui	$s0, 1
memory[265] <= 32'h00000000;	//			nop
memory[266] <= 32'h00000000;	//			nop
memory[267] <= 32'h00000000;	//			nop
memory[268] <= 32'h00000000;	//			nop
memory[269] <= 32'h00000000;	//			nop
memory[270] <= 32'h0601000b;	//			bgez	$s0, branch8
memory[271] <= 32'h00000000;	//			nop
memory[272] <= 32'h00000000;	//			nop
memory[273] <= 32'h00000000;	//			nop
memory[274] <= 32'h00000000;	//			nop
memory[275] <= 32'h00000000;	//			nop
memory[276] <= 32'h0800013e;	//			j	error
memory[277] <= 32'h00000000;	//			nop
memory[278] <= 32'h00000000;	//			nop
memory[279] <= 32'h00000000;	//			nop
memory[280] <= 32'h00000000;	//			nop
memory[281] <= 32'h00000000;	//			nop
memory[282] <= 32'h08000126;	//	branch8:	j	jump1
memory[283] <= 32'h00000000;	//			nop
memory[284] <= 32'h00000000;	//			nop
memory[285] <= 32'h00000000;	//			nop
memory[286] <= 32'h00000000;	//			nop
memory[287] <= 32'h00000000;	//			nop
memory[288] <= 32'h2210fffe;	//			addi	$s0, $s0, -2
memory[289] <= 32'h00000000;	//			nop
memory[290] <= 32'h00000000;	//			nop
memory[291] <= 32'h00000000;	//			nop
memory[292] <= 32'h00000000;	//			nop
memory[293] <= 32'h00000000;	//			nop
memory[294] <= 32'h0c000132;	//	jump1:		jal	jal1
memory[295] <= 32'h00000000;	//			nop
memory[296] <= 32'h00000000;	//			nop
memory[297] <= 32'h00000000;	//			nop
memory[298] <= 32'h00000000;	//			nop
memory[299] <= 32'h00000000;	//			nop
memory[300] <= 32'h08000018;	//			j	start
memory[301] <= 32'h00000000;	//			nop
memory[302] <= 32'h00000000;	//			nop
memory[303] <= 32'h00000000;	//			nop
memory[304] <= 32'h00000000;	//			nop
memory[305] <= 32'h00000000;	//			nop
memory[306] <= 32'h00000000;	//	jal1:		jr	$ra
memory[307] <= 32'h03e00008;	//			nop
memory[308] <= 32'h00000000;	//			nop
memory[309] <= 32'h00000000;	//			nop
memory[310] <= 32'h00000000;	//			nop
memory[311] <= 32'h00000000;	//			nop
memory[312] <= 32'h00000000;	//			j	error
memory[313] <= 32'h0800013e;	//			nop
memory[314] <= 32'h00000000;	//			nop
memory[315] <= 32'h00000000;	//			nop
memory[316] <= 32'h00000000;	//			nop
memory[317] <= 32'h00000000;	//			nop
memory[318] <= 32'h00000008;	//	error:		jr	$zero
memory[319] <= 32'h00000000;	//			nop
memory[320] <= 32'h00000000;	//			nop
memory[321] <= 32'h00000000;	//			nop
memory[322] <= 32'h00000000;	//			nop
memory[323] <= 32'h00000000;	//			nop
memory[324] <= 32'h00000000;	//			ori	$v0, $zero, 10
memory[325] <= 32'h3402000a;	//			nop
memory[326] <= 32'h00000000;	//			nop
memory[327] <= 32'h00000000;	//			nop
memory[328] <= 32'h00000000;	//			nop
memory[329] <= 32'h00000000;	//			nop
memory[330] <= 32'h00000000;	//			nop
memory[331] <= 32'h00000000;	//			nop
memory[332] <= 32'h00000000;	//			nop
memory[333] <= 32'h00000000;	//			nop
memory[334] <= 32'h00000000;	//			nop
memory[335] <= 32'h00000000;	//			nop
*/




/*
Memory[0] = 32'h34040000;
Memory[1] = 32'h00000000;
Memory[2] = 32'h00000000;
Memory[3] = 32'h00000000;
Memory[4] = 32'h00000000;
Memory[5] = 32'h00000000;
Memory[6] = 32'h08000018;
Memory[7] = 32'h00000000;
Memory[8] = 32'h00000000;
Memory[9] = 32'h00000000;
Memory[10] = 32'h00000000;
Memory[11] = 32'h00000000;
Memory[12] = 32'h2004000a;
Memory[13] = 32'h00000000;
Memory[14] = 32'h00000000;
Memory[15] = 32'h00000000;
Memory[16] = 32'h00000000;
Memory[17] = 32'h00000000;
Memory[18] = 32'h2004000a;
Memory[19] = 32'h00000000;
Memory[20] = 32'h00000000;
Memory[21] = 32'h00000000;
Memory[22] = 32'h00000000;
Memory[23] = 32'h00000000;
Memory[24] = 32'h8c900004;
Memory[25] = 32'h00000000;
Memory[26] = 32'h00000000;
Memory[27] = 32'h00000000;
Memory[28] = 32'h00000000;
Memory[29] = 32'h00000000;
Memory[30] = 32'h8c900008;
Memory[31] = 32'h00000000;
Memory[32] = 32'h00000000;
Memory[33] = 32'h00000000;
Memory[34] = 32'h00000000;
Memory[35] = 32'h00000000;
Memory[36] = 32'hac900000;
Memory[37] = 32'h00000000;
Memory[38] = 32'h00000000;
Memory[39] = 32'h00000000;
Memory[40] = 32'h00000000;
Memory[41] = 32'h00000000;
Memory[42] = 32'hac90000c;
Memory[43] = 32'h00000000;
Memory[44] = 32'h00000000;
Memory[45] = 32'h00000000;
Memory[46] = 32'h00000000;
Memory[47] = 32'h00000000;
Memory[48] = 32'h8c910000;
Memory[49] = 32'h00000000;
Memory[50] = 32'h00000000;
Memory[51] = 32'h00000000;
Memory[52] = 32'h00000000;
Memory[53] = 32'h00000000;
Memory[54] = 32'h8c92000c;
Memory[55] = 32'h00000000;
Memory[56] = 32'h00000000;
Memory[57] = 32'h00000000;
Memory[58] = 32'h00000000;
Memory[59] = 32'h00000000;
Memory[60] = 32'h12000017;
Memory[61] = 32'h00000000;
Memory[62] = 32'h00000000;
Memory[63] = 32'h00000000;
Memory[64] = 32'h00000000;
Memory[65] = 32'h00000000;
Memory[66] = 32'h02008820;
Memory[67] = 32'h00000000;
Memory[68] = 32'h00000000;
Memory[69] = 32'h00000000;
Memory[70] = 32'h00000000;
Memory[71] = 32'h00000000;
Memory[72] = 32'h1211000b;
Memory[73] = 32'h00000000;
Memory[74] = 32'h00000000;
Memory[75] = 32'h00000000;
Memory[76] = 32'h00000000;
Memory[77] = 32'h00000000;
Memory[78] = 32'h0800013e;
Memory[79] = 32'h00000000;
Memory[80] = 32'h00000000;
Memory[81] = 32'h00000000;
Memory[82] = 32'h00000000;
Memory[83] = 32'h00000000;
Memory[84] = 32'h2010ffff;
Memory[85] = 32'h00000000;
Memory[86] = 32'h00000000;
Memory[87] = 32'h00000000;
Memory[88] = 32'h00000000;
Memory[89] = 32'h00000000;
Memory[90] = 32'h0601ffbd;
Memory[91] = 32'h00000000;
Memory[92] = 32'h00000000;
Memory[93] = 32'h00000000;
Memory[94] = 32'h00000000;
Memory[95] = 32'h00000000;
Memory[96] = 32'h22100001;
Memory[97] = 32'h00000000;
Memory[98] = 32'h00000000;
Memory[99] = 32'h00000000;
Memory[100] = 32'h00000000;
Memory[101] = 32'h00000000;
Memory[102] = 32'h0601000b;
Memory[103] = 32'h00000000;
Memory[104] = 32'h00000000;
Memory[105] = 32'h00000000;
Memory[106] = 32'h00000000;
Memory[107] = 32'h00000000;
Memory[108] = 32'h0800013e;
Memory[109] = 32'h00000000;
Memory[110] = 32'h00000000;
Memory[111] = 32'h00000000;
Memory[112] = 32'h00000000;
Memory[113] = 32'h00000000;
Memory[114] = 32'h2010ffff;
Memory[115] = 32'h00000000;
Memory[116] = 32'h00000000;
Memory[117] = 32'h00000000;
Memory[118] = 32'h00000000;
Memory[119] = 32'h00000000;
Memory[120] = 32'h1e000017;
Memory[121] = 32'h00000000;
Memory[122] = 32'h00000000;
Memory[123] = 32'h00000000;
Memory[124] = 32'h00000000;
Memory[125] = 32'h00000000;
Memory[126] = 32'h20100001;
Memory[127] = 32'h00000000;
Memory[128] = 32'h00000000;
Memory[129] = 32'h00000000;
Memory[130] = 32'h00000000;
Memory[131] = 32'h00000000;
Memory[132] = 32'h1e00000b;
Memory[133] = 32'h00000000;
Memory[134] = 32'h00000000;
Memory[135] = 32'h00000000;
Memory[136] = 32'h00000000;
Memory[137] = 32'h00000000;
Memory[138] = 32'h0800013e;
Memory[139] = 32'h00000000;
Memory[140] = 32'h00000000;
Memory[141] = 32'h00000000;
Memory[142] = 32'h00000000;
Memory[143] = 32'h00000000;
Memory[144] = 32'h06000017;
Memory[145] = 32'h00000000;
Memory[146] = 32'h00000000;
Memory[147] = 32'h00000000;
Memory[148] = 32'h00000000;
Memory[149] = 32'h00000000;
Memory[150] = 32'h2010ffff;
Memory[151] = 32'h00000000;
Memory[152] = 32'h00000000;
Memory[153] = 32'h00000000;
Memory[154] = 32'h00000000;
Memory[155] = 32'h00000000;
Memory[156] = 32'h0600000b;
Memory[157] = 32'h00000000;
Memory[158] = 32'h00000000;
Memory[159] = 32'h00000000;
Memory[160] = 32'h00000000;
Memory[161] = 32'h00000000;
Memory[162] = 32'h0800013e;
Memory[163] = 32'h00000000;
Memory[164] = 32'h00000000;
Memory[165] = 32'h00000000;
Memory[166] = 32'h00000000;
Memory[167] = 32'h00000000;
Memory[168] = 32'h2011ffff;
Memory[169] = 32'h00000000;
Memory[170] = 32'h00000000;
Memory[171] = 32'h00000000;
Memory[172] = 32'h00000000;
Memory[173] = 32'h00000000;
Memory[174] = 32'h16110011;
Memory[175] = 32'h00000000;
Memory[176] = 32'h00000000;
Memory[177] = 32'h00000000;
Memory[178] = 32'h00000000;
Memory[179] = 32'h00000000;
Memory[180] = 32'h1600000b;
Memory[181] = 32'h00000000;
Memory[182] = 32'h00000000;
Memory[183] = 32'h00000000;
Memory[184] = 32'h00000000;
Memory[185] = 32'h00000000;
Memory[186] = 32'h0800013e;
Memory[187] = 32'h00000000;
Memory[188] = 32'h00000000;
Memory[189] = 32'h00000000;
Memory[190] = 32'h00000000;
Memory[191] = 32'h00000000;
Memory[192] = 32'h20100080;
Memory[193] = 32'h00000000;
Memory[194] = 32'h00000000;
Memory[195] = 32'h00000000;
Memory[196] = 32'h00000000;
Memory[197] = 32'h00000000;
Memory[198] = 32'ha0900000;
Memory[199] = 32'h00000000;
Memory[200] = 32'h00000000;
Memory[201] = 32'h00000000;
Memory[202] = 32'h00000000;
Memory[203] = 32'h00000000;
Memory[204] = 32'h80900000;
Memory[205] = 32'h00000000;
Memory[206] = 32'h00000000;
Memory[207] = 32'h00000000;
Memory[208] = 32'h00000000;
Memory[209] = 32'h00000000;
Memory[210] = 32'h1a00000b;
Memory[211] = 32'h00000000;
Memory[212] = 32'h00000000;
Memory[213] = 32'h00000000;
Memory[214] = 32'h00000000;
Memory[215] = 32'h00000000;
Memory[216] = 32'h0800013e;
Memory[217] = 32'h00000000;
Memory[218] = 32'h00000000;
Memory[219] = 32'h00000000;
Memory[220] = 32'h00000000;
Memory[221] = 32'h00000000;
Memory[222] = 32'h2010ffff;
Memory[223] = 32'h00000000;
Memory[224] = 32'h00000000;
Memory[225] = 32'h00000000;
Memory[226] = 32'h00000000;
Memory[227] = 32'h00000000;
Memory[228] = 32'ha4900000;
Memory[229] = 32'h00000000;
Memory[230] = 32'h00000000;
Memory[231] = 32'h00000000;
Memory[232] = 32'h00000000;
Memory[233] = 32'h00000000;
Memory[234] = 32'h20100000;
Memory[235] = 32'h00000000;
Memory[236] = 32'h00000000;
Memory[237] = 32'h00000000;
Memory[238] = 32'h00000000;
Memory[239] = 32'h00000000;
Memory[240] = 32'h84900000;
Memory[241] = 32'h00000000;
Memory[242] = 32'h00000000;
Memory[243] = 32'h00000000;
Memory[244] = 32'h00000000;
Memory[245] = 32'h00000000;
Memory[246] = 32'h1a00000b;
Memory[247] = 32'h00000000;
Memory[248] = 32'h00000000;
Memory[249] = 32'h00000000;
Memory[250] = 32'h00000000;
Memory[251] = 32'h00000000;
Memory[252] = 32'h0800013e;
Memory[253] = 32'h00000000;
Memory[254] = 32'h00000000;
Memory[255] = 32'h00000000;
Memory[256] = 32'h00000000;
Memory[257] = 32'h00000000;
Memory[258] = 32'h2010ffff;
Memory[259] = 32'h00000000;
Memory[260] = 32'h00000000;
Memory[261] = 32'h00000000;
Memory[262] = 32'h00000000;
Memory[263] = 32'h00000000;
Memory[264] = 32'h3c100001;
Memory[265] = 32'h00000000;
Memory[266] = 32'h00000000;
Memory[267] = 32'h00000000;
Memory[268] = 32'h00000000;
Memory[269] = 32'h00000000;
Memory[270] = 32'h0601000b;
Memory[271] = 32'h00000000;
Memory[272] = 32'h00000000;
Memory[273] = 32'h00000000;
Memory[274] = 32'h00000000;
Memory[275] = 32'h00000000;
Memory[276] = 32'h0800013e;
Memory[277] = 32'h00000000;
Memory[278] = 32'h00000000;
Memory[279] = 32'h00000000;
Memory[280] = 32'h00000000;
Memory[281] = 32'h00000000;
Memory[282] = 32'h08000126;
Memory[283] = 32'h00000000;
Memory[284] = 32'h00000000;
Memory[285] = 32'h00000000;
Memory[286] = 32'h00000000;
Memory[287] = 32'h00000000;
Memory[288] = 32'h2210fffe;
Memory[289] = 32'h00000000;
Memory[290] = 32'h00000000;
Memory[291] = 32'h00000000;
Memory[292] = 32'h00000000;
Memory[293] = 32'h00000000;
Memory[294] = 32'h0c000132;
Memory[295] = 32'h00000000;
Memory[296] = 32'h00000000;
Memory[297] = 32'h00000000;
Memory[298] = 32'h00000000;
Memory[299] = 32'h00000000;
Memory[300] = 32'h08000018;
Memory[301] = 32'h00000000;
Memory[302] = 32'h00000000;
Memory[303] = 32'h00000000;
Memory[304] = 32'h00000000;
Memory[305] = 32'h00000000;
Memory[306] = 32'h03e00008;
Memory[307] = 32'h00000000;
Memory[308] = 32'h00000000;
Memory[309] = 32'h00000000;
Memory[310] = 32'h00000000;
Memory[311] = 32'h00000000;
Memory[312] = 32'h0800013e;
Memory[313] = 32'h00000000;
Memory[314] = 32'h00000000;
Memory[315] = 32'h00000000;
Memory[316] = 32'h00000000;
Memory[317] = 32'h00000000;
Memory[318] = 32'h00000008;
Memory[319] = 32'h00000000;
Memory[320] = 32'h00000000;
Memory[321] = 32'h00000000;
Memory[322] = 32'h00000000;
Memory[323] = 32'h00000000;
Memory[324] = 32'h3402000a;
Memory[325] = 32'h00000000;
Memory[326] = 32'h00000000;
Memory[327] = 32'h00000000;
Memory[328] = 32'h00000000;
Memory[329] = 32'h00000000;
Memory[330] = 32'h00000000;
Memory[331] = 32'h00000000;
Memory[332] = 32'h00000000;
Memory[333] = 32'h00000000;
Memory[334] = 32'h00000000;
Memory[335] = 32'h00000000;
*/


/*
//          Public Test Case Labs 9-14 
    Memory[0] = 32'h20100001;
    Memory[1] = 32'h00000000;
    Memory[2] = 32'h00000000;
    Memory[3] = 32'h00000000;
    Memory[4] = 32'h00000000;
    Memory[5] = 32'h00000000;
    Memory[6] = 32'h20110001;
    Memory[7] = 32'h00000000;
    Memory[8] = 32'h00000000;
    Memory[9] = 32'h00000000;
    Memory[10] = 32'h00000000;
    Memory[11] = 32'h00000000;
    Memory[12] = 32'h02118024;
    Memory[13] = 32'h00000000;
    Memory[14] = 32'h00000000;
    Memory[15] = 32'h00000000;
    Memory[16] = 32'h00000000;
    Memory[17] = 32'h00000000;
    Memory[18] = 32'h02008024;
    Memory[19] = 32'h00000000;
    Memory[20] = 32'h00000000;
    Memory[21] = 32'h00000000;
    Memory[22] = 32'h00000000;
    Memory[23] = 32'h00000000;
    Memory[24] = 32'h02308022;
    Memory[25] = 32'h00000000;
    Memory[26] = 32'h00000000;
    Memory[27] = 32'h00000000;
    Memory[28] = 32'h00000000;
    Memory[29] = 32'h00000000;
    Memory[30] = 32'h02008027;
    Memory[31] = 32'h00000000;
    Memory[32] = 32'h00000000;
    Memory[33] = 32'h00000000;
    Memory[34] = 32'h00000000;
    Memory[35] = 32'h00000000;
    Memory[36] = 32'h02008027;
    Memory[37] = 32'h00000000;
    Memory[38] = 32'h00000000;
    Memory[39] = 32'h00000000;
    Memory[40] = 32'h00000000;
    Memory[41] = 32'h00000000;
    Memory[42] = 32'h00008025;
    Memory[43] = 32'h00000000;
    Memory[44] = 32'h00000000;
    Memory[45] = 32'h00000000;
    Memory[46] = 32'h00000000;
    Memory[47] = 32'h00000000;
    Memory[48] = 32'h02208025;
    Memory[49] = 32'h00000000;
    Memory[50] = 32'h00000000;
    Memory[51] = 32'h00000000;
    Memory[52] = 32'h00000000;
    Memory[53] = 32'h00000000;
    Memory[54] = 32'h00108080;
    Memory[55] = 32'h00000000;
    Memory[56] = 32'h00000000;
    Memory[57] = 32'h00000000;
    Memory[58] = 32'h00000000;
    Memory[59] = 32'h00000000;
    Memory[60] = 32'h02308004;
    Memory[61] = 32'h00000000;
    Memory[62] = 32'h00000000;
    Memory[63] = 32'h00000000;
    Memory[64] = 32'h00000000;
    Memory[65] = 32'h00000000;
    Memory[66] = 32'h0200802a;
    Memory[67] = 32'h00000000;
    Memory[68] = 32'h00000000;
    Memory[69] = 32'h00000000;
    Memory[70] = 32'h00000000;
    Memory[71] = 32'h00000000;
    Memory[72] = 32'h0211802a;
    Memory[73] = 32'h00000000;
    Memory[74] = 32'h00000000;
    Memory[75] = 32'h00000000;
    Memory[76] = 32'h00000000;
    Memory[77] = 32'h00000000;
    Memory[78] = 32'h00118043;
    Memory[79] = 32'h00000000;
    Memory[80] = 32'h00000000;
    Memory[81] = 32'h00000000;
    Memory[82] = 32'h00000000;
    Memory[83] = 32'h00000000;
    Memory[84] = 32'h00118007;
    Memory[85] = 32'h00000000;
    Memory[86] = 32'h00000000;
    Memory[87] = 32'h00000000;
    Memory[88] = 32'h00000000;
    Memory[89] = 32'h00000000;
    Memory[90] = 32'h00118042;
    Memory[91] = 32'h00000000;
    Memory[92] = 32'h00000000;
    Memory[93] = 32'h00000000;
    Memory[94] = 32'h00000000;
    Memory[95] = 32'h00000000;
    Memory[96] = 32'h001180c0;
    Memory[97] = 32'h00000000;
    Memory[98] = 32'h00000000;
    Memory[99] = 32'h00000000;
    Memory[100] = 32'h00000000;
    Memory[101] = 32'h00000000;
    Memory[102] = 32'h001080c2;
    Memory[103] = 32'h00000000;
    Memory[104] = 32'h00000000;
    Memory[105] = 32'h00000000;
    Memory[106] = 32'h00000000;
    Memory[107] = 32'h00000000;
    Memory[108] = 32'h02308004;
    Memory[109] = 32'h00000000;
    Memory[110] = 32'h00000000;
    Memory[111] = 32'h00000000;
    Memory[112] = 32'h00000000;
    Memory[113] = 32'h00000000;
    Memory[114] = 32'h02308006;
    Memory[115] = 32'h00000000;
    Memory[116] = 32'h00000000;
    Memory[117] = 32'h00000000;
    Memory[118] = 32'h00000000;
    Memory[119] = 32'h00000000;
    Memory[120] = 32'h02118026;
    Memory[121] = 32'h00000000;
    Memory[122] = 32'h00000000;
    Memory[123] = 32'h00000000;
    Memory[124] = 32'h00000000;
    Memory[125] = 32'h00000000;
    Memory[126] = 32'h02118026;
    Memory[127] = 32'h00000000;
    Memory[128] = 32'h00000000;
    Memory[129] = 32'h00000000;
    Memory[130] = 32'h00000000;
    Memory[131] = 32'h00000000;
    Memory[132] = 32'h20120004;
    Memory[133] = 32'h00000000;
    Memory[134] = 32'h00000000;
    Memory[135] = 32'h00000000;
    Memory[136] = 32'h00000000;
    Memory[137] = 32'h00000000;
    Memory[138] = 32'h72128002;
    Memory[139] = 32'h00000000;
    Memory[140] = 32'h00000000;
    Memory[141] = 32'h00000000;
    Memory[142] = 32'h00000000;
    Memory[143] = 32'h00000000;
    Memory[144] = 32'h22100004;
    Memory[145] = 32'h00000000;
    Memory[146] = 32'h00000000;
    Memory[147] = 32'h00000000;
    Memory[148] = 32'h00000000;
    Memory[149] = 32'h00000000;
    Memory[150] = 32'h32100000;
    Memory[151] = 32'h00000000;
    Memory[152] = 32'h00000000;
    Memory[153] = 32'h00000000;
    Memory[154] = 32'h00000000;
    Memory[155] = 32'h00000000;
    Memory[156] = 32'h36100001;
    Memory[157] = 32'h00000000;
    Memory[158] = 32'h00000000;
    Memory[159] = 32'h00000000;
    Memory[160] = 32'h00000000;
    Memory[161] = 32'h00000000;
    Memory[162] = 32'h2a100000;
    Memory[163] = 32'h00000000;
    Memory[164] = 32'h00000000;
    Memory[165] = 32'h00000000;
    Memory[166] = 32'h00000000;
    Memory[167] = 32'h00000000;
    Memory[168] = 32'h2a100001;
    Memory[169] = 32'h00000000;
    Memory[170] = 32'h00000000;
    Memory[171] = 32'h00000000;
    Memory[172] = 32'h00000000;
    Memory[173] = 32'h00000000;
    Memory[174] = 32'h3a100001;
    Memory[175] = 32'h00000000;
    Memory[176] = 32'h00000000;
    Memory[177] = 32'h00000000;
    Memory[178] = 32'h00000000;
    Memory[179] = 32'h00000000;
    Memory[180] = 32'h3a100001;
    Memory[181] = 32'h00000000;
    Memory[182] = 32'h00000000;
    Memory[183] = 32'h00000000;
    Memory[184] = 32'h00000000;
    Memory[185] = 32'h00000000;
    Memory[186] = 32'h2010fffe;
    Memory[187] = 32'h00000000;
    Memory[188] = 32'h00000000;
    Memory[189] = 32'h00000000;
    Memory[190] = 32'h00000000;
    Memory[191] = 32'h00000000;
    Memory[192] = 32'h20110002;
    Memory[193] = 32'h00000000;
    Memory[194] = 32'h00000000;
    Memory[195] = 32'h00000000;
    Memory[196] = 32'h00000000;
    Memory[197] = 32'h00000000;
    Memory[198] = 32'h0230902b;
    Memory[199] = 32'h00000000;
    Memory[200] = 32'h00000000;
    Memory[201] = 32'h00000000;
    Memory[202] = 32'h00000000;
    Memory[203] = 32'h00000000;
    Memory[204] = 32'h2e30fffe;
    Memory[205] = 32'h00000000;
    Memory[206] = 32'h00000000;
    Memory[207] = 32'h00000000;
    Memory[208] = 32'h00000000;
    Memory[209] = 32'h00000000;
    Memory[210] = 32'h0220800a;
    Memory[211] = 32'h00000000;
    Memory[212] = 32'h00000000;
    Memory[213] = 32'h00000000;
    Memory[214] = 32'h00000000;
    Memory[215] = 32'h00000000;
    Memory[216] = 32'h0011800b;
    Memory[217] = 32'h00000000;
    Memory[218] = 32'h00000000;
    Memory[219] = 32'h00000000;
    Memory[220] = 32'h00000000;
    Memory[221] = 32'h00000000;
    Memory[222] = 32'h02328020;
    Memory[223] = 32'h00000000;
    Memory[224] = 32'h00000000;
    Memory[225] = 32'h00000000;
    Memory[226] = 32'h00000000;
    Memory[227] = 32'h00000000;
    Memory[228] = 32'h2010fffe;
    Memory[229] = 32'h00000000;
    Memory[230] = 32'h00000000;
    Memory[231] = 32'h00000000;
    Memory[232] = 32'h00000000;
    Memory[233] = 32'h00000000;
    Memory[234] = 32'h02308821;
    Memory[235] = 32'h00000000;
    Memory[236] = 32'h00000000;
    Memory[237] = 32'h00000000;
    Memory[238] = 32'h00000000;
    Memory[239] = 32'h00000000;
    Memory[240] = 32'h2411ffff;
    Memory[241] = 32'h00000000;
    Memory[242] = 32'h00000000;
    Memory[243] = 32'h00000000;
    Memory[244] = 32'h00000000;
    Memory[245] = 32'h00000000;
    Memory[246] = 32'h20120020;
    Memory[247] = 32'h00000000;
    Memory[248] = 32'h00000000;
    Memory[249] = 32'h00000000;
    Memory[250] = 32'h00000000;
    Memory[251] = 32'h00000000;
    Memory[252] = 32'h02320018;
    Memory[253] = 32'h00000000;
    Memory[254] = 32'h00000000;
    Memory[255] = 32'h00000000;
    Memory[256] = 32'h00000000;
    Memory[257] = 32'h00000000;
    Memory[258] = 32'h0000a010;
    Memory[259] = 32'h00000000;
    Memory[260] = 32'h00000000;
    Memory[261] = 32'h00000000;
    Memory[262] = 32'h00000000;
    Memory[263] = 32'h00000000;
    Memory[264] = 32'h0000a812;
    Memory[265] = 32'h00000000;
    Memory[266] = 32'h00000000;
    Memory[267] = 32'h00000000;
    Memory[268] = 32'h00000000;
    Memory[269] = 32'h00000000;
    Memory[270] = 32'h02320019;
    Memory[271] = 32'h00000000;
    Memory[272] = 32'h00000000;
    Memory[273] = 32'h00000000;
    Memory[274] = 32'h00000000;
    Memory[275] = 32'h00000000;
    Memory[276] = 32'h0000a010;
    Memory[277] = 32'h00000000;
    Memory[278] = 32'h00000000;
    Memory[279] = 32'h00000000;
    Memory[280] = 32'h00000000;
    Memory[281] = 32'h00000000;
    Memory[282] = 32'h0000a812;
    Memory[283] = 32'h00000000;
    Memory[284] = 32'h00000000;
    Memory[285] = 32'h00000000;
    Memory[286] = 32'h00000000;
    Memory[287] = 32'h00000000;
    Memory[288] = 32'h72320000;
    Memory[289] = 32'h00000000;
    Memory[290] = 32'h00000000;
    Memory[291] = 32'h00000000;
    Memory[292] = 32'h00000000;
    Memory[293] = 32'h00000000;
    Memory[294] = 32'h0000a010;
    Memory[295] = 32'h00000000;
    Memory[296] = 32'h00000000;
    Memory[297] = 32'h00000000;
    Memory[298] = 32'h00000000;
    Memory[299] = 32'h00000000;
    Memory[300] = 32'h0000a812;
    Memory[301] = 32'h00000000;
    Memory[302] = 32'h00000000;
    Memory[303] = 32'h00000000;
    Memory[304] = 32'h00000000;
    Memory[305] = 32'h00000000;
    Memory[306] = 32'h02400011;
    Memory[307] = 32'h00000000;
    Memory[308] = 32'h00000000;
    Memory[309] = 32'h00000000;
    Memory[310] = 32'h00000000;
    Memory[311] = 32'h00000000;
    Memory[312] = 32'h02200013;
    Memory[313] = 32'h00000000;
    Memory[314] = 32'h00000000;
    Memory[315] = 32'h00000000;
    Memory[316] = 32'h00000000;
    Memory[317] = 32'h00000000;
    Memory[318] = 32'h0000a010;
    Memory[319] = 32'h00000000;
    Memory[320] = 32'h00000000;
    Memory[321] = 32'h00000000;
    Memory[322] = 32'h00000000;
    Memory[323] = 32'h00000000;
    Memory[324] = 32'h0000a812;
    Memory[325] = 32'h00000000;
    Memory[326] = 32'h00000000;
    Memory[327] = 32'h00000000;
    Memory[328] = 32'h00000000;
    Memory[329] = 32'h00000000;
    Memory[330] = 32'h3231ffff;
    Memory[331] = 32'h00000000;
    Memory[332] = 32'h00000000;
    Memory[333] = 32'h00000000;
    Memory[334] = 32'h00000000;
    Memory[335] = 32'h00000000;
    Memory[336] = 32'h72920004;
    Memory[337] = 32'h00000000;
    Memory[338] = 32'h00000000;
    Memory[339] = 32'h00000000;
    Memory[340] = 32'h00000000;
    Memory[341] = 32'h00000000;
    Memory[342] = 32'h0000a010;
    Memory[343] = 32'h00000000;
    Memory[344] = 32'h00000000;
    Memory[345] = 32'h00000000;
    Memory[346] = 32'h00000000;
    Memory[347] = 32'h00000000;
    Memory[348] = 32'h0000a812;
    Memory[349] = 32'h00000000;
    Memory[350] = 32'h00000000;
    Memory[351] = 32'h00000000;
    Memory[352] = 32'h00000000;
    Memory[353] = 32'h00000000;
    Memory[354] = 32'h20120001;
    Memory[355] = 32'h00000000;
    Memory[356] = 32'h00000000;
    Memory[357] = 32'h00000000;
    Memory[358] = 32'h00000000;
    Memory[359] = 32'h00000000;
    Memory[360] = 32'h00328fc2;
    Memory[361] = 32'h00000000;
    Memory[362] = 32'h00000000;
    Memory[363] = 32'h00000000;
    Memory[364] = 32'h00000000;
    Memory[365] = 32'h00000000;
    Memory[366] = 32'h2014001f;
    Memory[367] = 32'h00000000;
    Memory[368] = 32'h00000000;
    Memory[369] = 32'h00000000;
    Memory[370] = 32'h00000000;
    Memory[371] = 32'h00000000;
    Memory[372] = 32'h02918846;
    Memory[373] = 32'h00000000;
    Memory[374] = 32'h00000000;
    Memory[375] = 32'h00000000;
    Memory[376] = 32'h00000000;
    Memory[377] = 32'h00000000;
    Memory[378] = 32'h34110FF0;
    Memory[379] = 32'h00000000;
    Memory[380] = 32'h00000000;
    Memory[381] = 32'h00000000;
    Memory[382] = 32'h00000000;
    Memory[383] = 32'h00000000;
    Memory[384] = 32'h7c11a420;
    Memory[385] = 32'h00000000;
    Memory[386] = 32'h00000000;
    Memory[387] = 32'h00000000;
    Memory[388] = 32'h00000000;
    Memory[389] = 32'h00000000;
    Memory[390] = 32'h7c11a620;
    Memory[391] = 32'h00000000;
    Memory[392] = 32'h00000000;
    Memory[393] = 32'h00000000;
    Memory[394] = 32'h00000000;
    Memory[395] = 32'h00000000;
*/






        /* Count up by 3's
        for (index = 0; index < 128; index = index + 1) begin
            Memory[index] = index * 3;
        end
        */
    end
    
    
    always @ Address begin
        Instruction = memory[Address[11:2]];
    end
    
    
endmodule
